module gw_gao(
    \pwm_cnt[18] ,
    \pwm_cnt[17] ,
    \pwm_cnt[16] ,
    \pwm_cnt[15] ,
    \pwm_cnt[14] ,
    \pwm_cnt[13] ,
    \pwm_cnt[12] ,
    \pwm_cnt[11] ,
    \pwm_cnt[10] ,
    \pwm_cnt[9] ,
    \pwm_cnt[8] ,
    \pwm_cnt[7] ,
    \pwm_cnt[6] ,
    \pwm_cnt[5] ,
    \pwm_cnt[4] ,
    \pwm_cnt[3] ,
    \pwm_cnt[2] ,
    \pwm_cnt[1] ,
    \pwm_cnt[0] ,
    \pwm_out2_u0/val_max[19] ,
    \pwm_out2_u0/val_max[18] ,
    \pwm_out2_u0/val_max[17] ,
    \pwm_out2_u0/val_max[16] ,
    \pwm_out2_u0/val_max[15] ,
    \pwm_out2_u0/val_max[14] ,
    \pwm_out2_u0/val_max[13] ,
    \pwm_out2_u0/val_max[12] ,
    \pwm_out2_u0/val_max[11] ,
    \pwm_out2_u0/val_max[10] ,
    \pwm_out2_u0/val_max[9] ,
    \pwm_out2_u0/val_max[8] ,
    \pwm_out2_u0/val_max[7] ,
    \pwm_out2_u0/val_max[6] ,
    \pwm_out2_u0/val_max[5] ,
    \pwm_out2_u0/val_max[4] ,
    \pwm_out2_u0/val_max[3] ,
    \pwm_out2_u0/val_max[2] ,
    \pwm_out2_u0/val_max[1] ,
    \pwm_out2_u0/val_max[0] ,
    \pwm_out2_u0/pwm_find[18] ,
    \pwm_out2_u0/pwm_find[17] ,
    \pwm_out2_u0/pwm_find[16] ,
    \pwm_out2_u0/pwm_find[15] ,
    \pwm_out2_u0/pwm_find[14] ,
    \pwm_out2_u0/pwm_find[13] ,
    \pwm_out2_u0/pwm_find[12] ,
    \pwm_out2_u0/pwm_find[11] ,
    \pwm_out2_u0/pwm_find[10] ,
    \pwm_out2_u0/pwm_find[9] ,
    \pwm_out2_u0/pwm_find[8] ,
    \pwm_out2_u0/pwm_find[7] ,
    \pwm_out2_u0/pwm_find[6] ,
    \pwm_out2_u0/pwm_find[5] ,
    \pwm_out2_u0/pwm_find[4] ,
    \pwm_out2_u0/pwm_find[3] ,
    \pwm_out2_u0/pwm_find[2] ,
    \pwm_out2_u0/pwm_find[1] ,
    \pwm_out2_u0/pwm_find[0] ,
    \px[10] ,
    \px[9] ,
    \px[8] ,
    \px[7] ,
    \px[6] ,
    \px[5] ,
    \px[4] ,
    \px[3] ,
    \px[2] ,
    \px[1] ,
    \px[0] ,
    \img_processor_u0/vga_mark_out_top_u0/py[10] ,
    \img_processor_u0/vga_mark_out_top_u0/py[9] ,
    \img_processor_u0/vga_mark_out_top_u0/py[8] ,
    \img_processor_u0/vga_mark_out_top_u0/py[7] ,
    \img_processor_u0/vga_mark_out_top_u0/py[6] ,
    \img_processor_u0/vga_mark_out_top_u0/py[5] ,
    \img_processor_u0/vga_mark_out_top_u0/py[4] ,
    \img_processor_u0/vga_mark_out_top_u0/py[3] ,
    \img_processor_u0/vga_mark_out_top_u0/py[2] ,
    \img_processor_u0/vga_mark_out_top_u0/py[1] ,
    \img_processor_u0/vga_mark_out_top_u0/py[0] ,
    I_rst_n,
    I_clk_50m,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \pwm_cnt[18] ;
input \pwm_cnt[17] ;
input \pwm_cnt[16] ;
input \pwm_cnt[15] ;
input \pwm_cnt[14] ;
input \pwm_cnt[13] ;
input \pwm_cnt[12] ;
input \pwm_cnt[11] ;
input \pwm_cnt[10] ;
input \pwm_cnt[9] ;
input \pwm_cnt[8] ;
input \pwm_cnt[7] ;
input \pwm_cnt[6] ;
input \pwm_cnt[5] ;
input \pwm_cnt[4] ;
input \pwm_cnt[3] ;
input \pwm_cnt[2] ;
input \pwm_cnt[1] ;
input \pwm_cnt[0] ;
input \pwm_out2_u0/val_max[19] ;
input \pwm_out2_u0/val_max[18] ;
input \pwm_out2_u0/val_max[17] ;
input \pwm_out2_u0/val_max[16] ;
input \pwm_out2_u0/val_max[15] ;
input \pwm_out2_u0/val_max[14] ;
input \pwm_out2_u0/val_max[13] ;
input \pwm_out2_u0/val_max[12] ;
input \pwm_out2_u0/val_max[11] ;
input \pwm_out2_u0/val_max[10] ;
input \pwm_out2_u0/val_max[9] ;
input \pwm_out2_u0/val_max[8] ;
input \pwm_out2_u0/val_max[7] ;
input \pwm_out2_u0/val_max[6] ;
input \pwm_out2_u0/val_max[5] ;
input \pwm_out2_u0/val_max[4] ;
input \pwm_out2_u0/val_max[3] ;
input \pwm_out2_u0/val_max[2] ;
input \pwm_out2_u0/val_max[1] ;
input \pwm_out2_u0/val_max[0] ;
input \pwm_out2_u0/pwm_find[18] ;
input \pwm_out2_u0/pwm_find[17] ;
input \pwm_out2_u0/pwm_find[16] ;
input \pwm_out2_u0/pwm_find[15] ;
input \pwm_out2_u0/pwm_find[14] ;
input \pwm_out2_u0/pwm_find[13] ;
input \pwm_out2_u0/pwm_find[12] ;
input \pwm_out2_u0/pwm_find[11] ;
input \pwm_out2_u0/pwm_find[10] ;
input \pwm_out2_u0/pwm_find[9] ;
input \pwm_out2_u0/pwm_find[8] ;
input \pwm_out2_u0/pwm_find[7] ;
input \pwm_out2_u0/pwm_find[6] ;
input \pwm_out2_u0/pwm_find[5] ;
input \pwm_out2_u0/pwm_find[4] ;
input \pwm_out2_u0/pwm_find[3] ;
input \pwm_out2_u0/pwm_find[2] ;
input \pwm_out2_u0/pwm_find[1] ;
input \pwm_out2_u0/pwm_find[0] ;
input \px[10] ;
input \px[9] ;
input \px[8] ;
input \px[7] ;
input \px[6] ;
input \px[5] ;
input \px[4] ;
input \px[3] ;
input \px[2] ;
input \px[1] ;
input \px[0] ;
input \img_processor_u0/vga_mark_out_top_u0/py[10] ;
input \img_processor_u0/vga_mark_out_top_u0/py[9] ;
input \img_processor_u0/vga_mark_out_top_u0/py[8] ;
input \img_processor_u0/vga_mark_out_top_u0/py[7] ;
input \img_processor_u0/vga_mark_out_top_u0/py[6] ;
input \img_processor_u0/vga_mark_out_top_u0/py[5] ;
input \img_processor_u0/vga_mark_out_top_u0/py[4] ;
input \img_processor_u0/vga_mark_out_top_u0/py[3] ;
input \img_processor_u0/vga_mark_out_top_u0/py[2] ;
input \img_processor_u0/vga_mark_out_top_u0/py[1] ;
input \img_processor_u0/vga_mark_out_top_u0/py[0] ;
input I_rst_n;
input I_clk_50m;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \pwm_cnt[18] ;
wire \pwm_cnt[17] ;
wire \pwm_cnt[16] ;
wire \pwm_cnt[15] ;
wire \pwm_cnt[14] ;
wire \pwm_cnt[13] ;
wire \pwm_cnt[12] ;
wire \pwm_cnt[11] ;
wire \pwm_cnt[10] ;
wire \pwm_cnt[9] ;
wire \pwm_cnt[8] ;
wire \pwm_cnt[7] ;
wire \pwm_cnt[6] ;
wire \pwm_cnt[5] ;
wire \pwm_cnt[4] ;
wire \pwm_cnt[3] ;
wire \pwm_cnt[2] ;
wire \pwm_cnt[1] ;
wire \pwm_cnt[0] ;
wire \pwm_out2_u0/val_max[19] ;
wire \pwm_out2_u0/val_max[18] ;
wire \pwm_out2_u0/val_max[17] ;
wire \pwm_out2_u0/val_max[16] ;
wire \pwm_out2_u0/val_max[15] ;
wire \pwm_out2_u0/val_max[14] ;
wire \pwm_out2_u0/val_max[13] ;
wire \pwm_out2_u0/val_max[12] ;
wire \pwm_out2_u0/val_max[11] ;
wire \pwm_out2_u0/val_max[10] ;
wire \pwm_out2_u0/val_max[9] ;
wire \pwm_out2_u0/val_max[8] ;
wire \pwm_out2_u0/val_max[7] ;
wire \pwm_out2_u0/val_max[6] ;
wire \pwm_out2_u0/val_max[5] ;
wire \pwm_out2_u0/val_max[4] ;
wire \pwm_out2_u0/val_max[3] ;
wire \pwm_out2_u0/val_max[2] ;
wire \pwm_out2_u0/val_max[1] ;
wire \pwm_out2_u0/val_max[0] ;
wire \pwm_out2_u0/pwm_find[18] ;
wire \pwm_out2_u0/pwm_find[17] ;
wire \pwm_out2_u0/pwm_find[16] ;
wire \pwm_out2_u0/pwm_find[15] ;
wire \pwm_out2_u0/pwm_find[14] ;
wire \pwm_out2_u0/pwm_find[13] ;
wire \pwm_out2_u0/pwm_find[12] ;
wire \pwm_out2_u0/pwm_find[11] ;
wire \pwm_out2_u0/pwm_find[10] ;
wire \pwm_out2_u0/pwm_find[9] ;
wire \pwm_out2_u0/pwm_find[8] ;
wire \pwm_out2_u0/pwm_find[7] ;
wire \pwm_out2_u0/pwm_find[6] ;
wire \pwm_out2_u0/pwm_find[5] ;
wire \pwm_out2_u0/pwm_find[4] ;
wire \pwm_out2_u0/pwm_find[3] ;
wire \pwm_out2_u0/pwm_find[2] ;
wire \pwm_out2_u0/pwm_find[1] ;
wire \pwm_out2_u0/pwm_find[0] ;
wire \px[10] ;
wire \px[9] ;
wire \px[8] ;
wire \px[7] ;
wire \px[6] ;
wire \px[5] ;
wire \px[4] ;
wire \px[3] ;
wire \px[2] ;
wire \px[1] ;
wire \px[0] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[10] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[9] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[8] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[7] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[6] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[5] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[4] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[3] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[2] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[1] ;
wire \img_processor_u0/vga_mark_out_top_u0/py[0] ;
wire I_rst_n;
wire I_clk_50m;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i(I_rst_n),
    .data_i({\pwm_cnt[18] ,\pwm_cnt[17] ,\pwm_cnt[16] ,\pwm_cnt[15] ,\pwm_cnt[14] ,\pwm_cnt[13] ,\pwm_cnt[12] ,\pwm_cnt[11] ,\pwm_cnt[10] ,\pwm_cnt[9] ,\pwm_cnt[8] ,\pwm_cnt[7] ,\pwm_cnt[6] ,\pwm_cnt[5] ,\pwm_cnt[4] ,\pwm_cnt[3] ,\pwm_cnt[2] ,\pwm_cnt[1] ,\pwm_cnt[0] ,\pwm_out2_u0/val_max[19] ,\pwm_out2_u0/val_max[18] ,\pwm_out2_u0/val_max[17] ,\pwm_out2_u0/val_max[16] ,\pwm_out2_u0/val_max[15] ,\pwm_out2_u0/val_max[14] ,\pwm_out2_u0/val_max[13] ,\pwm_out2_u0/val_max[12] ,\pwm_out2_u0/val_max[11] ,\pwm_out2_u0/val_max[10] ,\pwm_out2_u0/val_max[9] ,\pwm_out2_u0/val_max[8] ,\pwm_out2_u0/val_max[7] ,\pwm_out2_u0/val_max[6] ,\pwm_out2_u0/val_max[5] ,\pwm_out2_u0/val_max[4] ,\pwm_out2_u0/val_max[3] ,\pwm_out2_u0/val_max[2] ,\pwm_out2_u0/val_max[1] ,\pwm_out2_u0/val_max[0] ,\pwm_out2_u0/pwm_find[18] ,\pwm_out2_u0/pwm_find[17] ,\pwm_out2_u0/pwm_find[16] ,\pwm_out2_u0/pwm_find[15] ,\pwm_out2_u0/pwm_find[14] ,\pwm_out2_u0/pwm_find[13] ,\pwm_out2_u0/pwm_find[12] ,\pwm_out2_u0/pwm_find[11] ,\pwm_out2_u0/pwm_find[10] ,\pwm_out2_u0/pwm_find[9] ,\pwm_out2_u0/pwm_find[8] ,\pwm_out2_u0/pwm_find[7] ,\pwm_out2_u0/pwm_find[6] ,\pwm_out2_u0/pwm_find[5] ,\pwm_out2_u0/pwm_find[4] ,\pwm_out2_u0/pwm_find[3] ,\pwm_out2_u0/pwm_find[2] ,\pwm_out2_u0/pwm_find[1] ,\pwm_out2_u0/pwm_find[0] ,\px[10] ,\px[9] ,\px[8] ,\px[7] ,\px[6] ,\px[5] ,\px[4] ,\px[3] ,\px[2] ,\px[1] ,\px[0] ,\img_processor_u0/vga_mark_out_top_u0/py[10] ,\img_processor_u0/vga_mark_out_top_u0/py[9] ,\img_processor_u0/vga_mark_out_top_u0/py[8] ,\img_processor_u0/vga_mark_out_top_u0/py[7] ,\img_processor_u0/vga_mark_out_top_u0/py[6] ,\img_processor_u0/vga_mark_out_top_u0/py[5] ,\img_processor_u0/vga_mark_out_top_u0/py[4] ,\img_processor_u0/vga_mark_out_top_u0/py[3] ,\img_processor_u0/vga_mark_out_top_u0/py[2] ,\img_processor_u0/vga_mark_out_top_u0/py[1] ,\img_processor_u0/vga_mark_out_top_u0/py[0] }),
    .clk_i(I_clk_50m)
);

endmodule
//
// Written by Synplify Pro 
// Product Version "P-2019.03G-Beta4"
// Program "Synplify Pro", Mapper "mapgw, Build 1429R"
// Sun Nov 17 13:24:49 2019
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\e:\gowin_projects\myproj\myproj_blue2\temp\gao\ao_control\gw_con_parameter.v "
// file 6 "\e:\gowin_projects\myproj\myproj_blue2\temp\gao\ao_control\gw_con_top_define.v "
// file 7 "\e:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_con\gw_con_top.v "
// file 8 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
nGQjNTRggZWOT6sWc6oyraDUFLfWAO/HbLF6wXbCqXPNp9WCDJpv1rHVczOIVgncR/b0+UeSwebZ
OxlPzCeuO1qPl8FPTKiUyycPd+J0aSTr5vl+//g43DlAnrAZWpp+9NwkyX7Tl4KQV38q+/ZFnqAd
fKrxDpwkhDu4v9GmdKTtVryneeZJtk+qfqQLeux8ui4DI7WokBCiLCcnunBZc7zPDJ4RNHhhj/d6
kphLiA+2e7BZhQi3+S17OFvZZeAZqB9QHyWn8tsgCw/p96pTPtatJ/h1TGMYgxgbBmCeWweLMmye
bCwg5pbhghYptD2zVIQFJWuiylXMfypQ3ZpFdA==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
x5gHfLwQ9h6IkqXYFQsKYOoMTbgAOviKZwc0Vf339pYT772gCzJCT3UDF+YsUsYbK+Pq7BKRT6Uf
HBulNYuf7y+Ku9k8h5gb4vT0dUa4DG8OSdHb7R0AC/h0AeBTlns2hBJ4OSQGxyyNBp2s9HonSdOM
8ZWZFAphVVtPxikUpfU8q9qzyHTb9jMLF3VfqHt1hy3qcsmu5t+UPmv9c2zjTl4NXRMUl5483dXo
fMq4baFS/ju/wiHFuRhteazMg0mM6BfGhtM2aDlFaVzlnFbwItgar6Mu4Fk1u80ynR+wqXfj4ur2
96zU62Pm3UBbG8dYUGOAgfAhYDkhAs6USGbytQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7104)
`pragma protect data_block
S64wz9lq30aLaC+kL/X10osfDUSymmrQf6hdQCYuLnmlW6w0Fzin4aO0g/WUobnGsoCOY7+vwaK7
shINCGen4o92p7HrSWBdN+5Baowett5dwKHQqJmKXDf8kRu2EUM6L5usvI7gmjwb0Oqr0AOxGdMA
IEt240OIHMHC5+4DWcK1R5uW4oisAZTZ0NJomTQDaMYTf0vbCXRvBfHpZ4l5DtYYykQ+1wrCdaX8
sSH+7Kja8QmLHvKxnpa8f5JIgVG/ucAiaLjJCwWMxb9Jgg651lo4it+/5Tpuo5y2qsnz4H1JMNUn
Uj2Wb4mlOEYAAuxfOQgISpA8CPBcEc7sbHGRaiqACMoKpmzuzNxNUD8P5cv6ovUqQfJUioqy8RZU
ncsdMPHyh5mNATv+rgnC5o/KV93EFFByE293XvqXEYEjt9+B0tjML3MngPfTex/cJ2bRYI1Y29hm
XTL62PjJKbMzmK9NpFeIkHzsZDbc2u2z/BIavl6tVtDLm+SAcnppavWyK/5wQreqZ2yB53u9z2o8
LprLjQ9sr4VB4syjJwQmDoIF3R2IbM/QcfbvefBq4dq5wIAzfUOIsG7ArZLpKq5bpD2Zb8A9OHiX
uvKXXGCAt2zRRcVLod4NupUa6X2EHnU26zdjJmoMtd40HPn4cS1oNYsj8oDgnMRuf/Usf2EPCPzZ
zBwI1jWvbx/LDqAKeiJy5p6Z3ppYHfexLl4KVFJwvZN/UAIWIEdE4gMnasijR0V/X7zNIff2Z+mg
Vst3itLdrWLhIpU72gmh+FTfXmgP5G0QzeUXu+8N1eSeRol7/A0ii/TmT6olTEgp5qz99PEILD9D
dwbTqx6rbR/vbvZYn5A6MKVaJHf1Cf2AGsVHwSde1kyO3hEKtQ4r9nRWUIdDLZuN0jDbKAOGjSOj
cKQrNjYtn3fCdAE+vAydqBHJo0aNdCmOVR4Q2pRU6nYrm/btQlG2q7hLFtC/KPp2DUkDmxN8r+5B
jtXBUi4kv0tFiBkb0PSxuTRWBbmxgMHvu2TByRH6BUq6yGS45JSdbjpP0iYwguTga9uQlQJseJvN
j15bPLNnu23qzXFj4YABLhVMn3u2NXCFJtuYMqFQMW1J4orX1gR/oDz9x64hSD6+sdyOMqp9gEDe
0WZRRJAd6GzrepdeVLDl8wkUL5q2LruU+iqjEWV6S9w6E/+nxR01/BtxYLYurB06WOIux2dQ288m
+GGE3sZDqGx+4Z8RhX1zXr+jWRREuhScq0o8HakXzrQJ5d6LY3XsmvevNbnVF62XHGOq0jtREcXU
H1rGoR5lC3ijAvpx7b8Nk6N9VmI+ia0y17PcS32wivatHlatOvDz21513YSpkq/Yw2A6uJRl8KVH
Jj+kLgnAtJuMsFxxnHHDEd0DwbhpHYNlklIcez4hcNHHcW8UY+129G8pPPfxT0aJwrvc8xdF3FO5
zGC7rZuAhq3x1cJ/zlTFsepDtjwvqoqUCODzgXBkdDzWftJn68ittbbm+zbQzXZHy39+5j/0bQGq
xrYRoc7uHFk9KdSbpbDJdvad2clSy0ty9w4csPYjbsz+kkb94vouUIdy2WpnMkdbST/cPwsGLpfj
udJD5z0gsk2qDLqeePnl3U/C9moYz+Cw5pa2tiYU0V8BmX7+oShtCNHaGx/694KY617H2GQzy3oA
m7axRdZFb0Wf5dz0Nx2TmDvYGlw8284EwrgIzrOmqP0aBAPXESpUujnN+olGWShGRd5EtgOyQLgI
HhCppZtOjMPSKULg1NinMUMFPFZIn3dNlRGv2wFaiFFWDgFJnKxRNHujBhtdwAf3yifrXHjvjlq+
rdBW/36IfXTsD2Hk9yW8sCyFEJ8thBI9kX8v9IynnWfRY77pExP+MXu6n1mMsAGI5+NMIIvtD3/I
8xOHQ4Fm3nw61qa/ENEbZE2xLwnNBdbKhRkOJ5E61hofSr+tdUO7JXbd6HEDKhyQgNHJRVAlCaZg
nxVNBSyNe05LUxwkXsArTwvBn8XteTvnwreP7Rvd46oUPX9at5gkj45CfbJkoid5ejxoP7oRA8pc
b+LtAJCrMLquvMjrcRKEjqw+yyUwIcTu2KqmtaORXZbFfDMTQidCAL5iiZiQBMmtRO3/2JWSeO/z
yisWQmRAJxgLaoyfQTxLqqv183VR0dQI10GRQNDUNkuSEADQyOOj93ejJfRl7bMQft7oV6nVSCuQ
y4cjRGk4zWKW0i3x9RhGpv3MBr3PSrgrf0dmtM+SQAyshs8XMHzJevWf/0Y+78vbIDJJg1KwCgc5
uDOLVwDKf4yKpJU7loF9aKfWzRojoC/RpzyT9A68n5qc+QDWvPhUBWhrKN8weI5h0z8dGcwY+9z9
yED1Ockg4xGHaqcWGGWbPa5C1rZUCPgFkHsmyLX8W66yGl24nohnk0O/GNwCNhNzhVwQwtkawho2
o4AiWfYhdFKXouZ/racJoqYuoAV/t9cIMNZEG2q8vvHIXNf6/NB3QDyyNrxBmJYSwEABPH7rCvDI
rDzMLY7dGRZ1CgyuP2Ge2RY28vqO1sN05e4EbXxxz2GQTnvAf62+oTQg4B3cMKNkFUzO4xLyV4M4
A3r8mmGj/Kw5MHLbs8dl44f+P9vU/+N7IiQWRgPdfhrNIPYmrRRw0o3UEl5GQMa7ersm2H20+i3Y
FLw9medsYw903pVmzIBH2R1YUdNrYOquqVdI3cEjOHbVLruEmC9CEP6s8mRyi9ixwNK1ZGF7StYb
lYUvkpMh/FbEOutMh2dAYwuCQaKcUtQmP3d/SMDOgrDKXiJKqE6tzq7W5TDy5HWT/Y43/TdUF8BK
0jJX/krAu+lIqq+KfAkrBVy1aZR7TVrpuJptvSWUogS/ZKOQecBI+DScbiM3p7ZHod5X9Hlt+on0
Eix/WyX6Xh7Qr5AqZcNwvF6rTmcIBKjZv6j+y2Flnb7VMqDsTB8bAOoBRPnWW7yEWyy4GXrxoX8F
Pj4hlK/sGSmfTI1ioE/HOfBGFUrMTCaxpq3uOcMxBQeeNoZJzL1HfxDFntp0z1s/Rv/KJcGluUaU
LRAaH/I5r9XgOinwSRcjpBrxjS+uiwZXJu1JuCQz+pQcsbsP1hc1ZM12XHKr/G9/xkPgzCiMVkLk
E0wlaFyCxuwgxb889oZCDYq+huWYcNbgMGyi0aW+QYuE8Ha9YlNJf3A3XJxk8tTaxhWqXNp4THVn
ZU7UM9mZwAvK6ef4+/UugG5R0gLQMPPSa4+TeXQDgSYeCOWKs8fwhKrEpzgFgoPv1e20fd7MS/bU
Op1AIbsXYQcxcPvkx9+QPszLjD2V5z1vmt91ndI0sgzflNwbUVdkhMwrBYowMnJKdCru7q6mqi/a
mCV3l5rBjDVHh0LiICc4jMrrSo6EiLhNwWFJWowZWTCkUNIZNUKegYjpBs7gmpuwndeGNxVfXCZn
iVlTRNTIfWj2fb8GIQ/mJDa7hzFxv/21KhESvnTDuaEjy9HaxR0+OljsYi6owDKtW/cj4ei5Khnn
kKXigqdMoPQnBBy5+Dlu8xs2AWSIQa1wUyoGqjBATErO6LXslghIbgq3y3ExZTY5kf7IKKLBmQaz
YxJh3X/LJLQkgk7ePJveOrVRNEA1BMm4TdqAFj4pBlAUeMcilNPhQ+gX38QGT480Pc2RFSWW1+ZN
oefjAnTTwBcZ8z5Yac/0qMttIH0mDph96GRuSx8VEpQ0hr5VAkTVoUohABBRUHcb9Ls90mRafwUA
lbI3mwbhRsCkcsDJB4jutp3wOCt0BVnc3b2+PBN7AjQRSASl93ofLhAxfVQ03l1nSibvSWe1+wbG
2dUJy5u2M55OD1N5tEIcI6o95cLbNOx36bQSpDSigg8keHtqgKYe+fFnQZUWWXohOI5mATn5hRPV
KiZfXbB31Oa5A3DDm+jb5C4+D6mSI2LLcQZe6yknElDChlD9GQhlBTqUAG8cGVwlMftOZ5E8BwPe
rkBZP4Ih+w5WxPnkeYmydhqWLnoSSI6HIFK+gkJzsuTlBOU93wYBBG6Umg67l3bAjI4Xib3N5jiB
ZbFxokxItCnNtf1FFaLK0+2KHPTAPbuhOE2o2IYQpnab8Zegs05TYPyRSf2/7WpTtkDdiF7ejKlc
sPA+xM8N6R6Yrwakae3dS+Mu2Y6OntbT4U51BJmslkUEf0mWTY96RF1BVKUL5SVRgCqHRAeMyHaz
qHvSApD1czKbgf4i6g3q68umeUXAJJLiegmNd+yLjbdIGrlofjvBhlw3n6umwbU2Sqxw0NQM8HQ5
K6XxvdnDQ1OBfko4XHIFhhkhse8agYli7HJ0cpOsC0vaeHoA+BTC0lAKOkOLLD9Q+wI5y2lOBRUI
R/+2kC8ndhlEWoROS1M+bMQ8AURisonhvfmHAt62wu6CSGlbYwkp1I3sUxtx9kMmPnGSe5NHe1Jr
wGSchJ1g/D0weviUf/8UAtojoJiQUi/eezHzww2DQfz5PvREUkVQC1Se72W8wF2L4ATqFFaua12b
wGFTzC1JLsaMMaPmL8v5S0d4vhhorHtY4uzrMjEeS8uzcjyssxaVOE/ZLklT7bX8DKdlmIhWRAKV
qHHvdKv7weZ9yTsxXKWZaUpg4MHP0v0gdGecJ8xkSageBrXGZp1pI47y6W0v7bc3EMyt7rV7D2nM
hwUGuqQhktdwoQiLapiHCtuLi1cKGeScbabmqW0gFXV5ooMTafetu2mHFAhx6q02YZAPQhfcosP/
gwCqIcK1YPBEyJ60SkW9/KGp/K4XCOuyqgbcI4RHUPXCHgI8cVy2pRTbCRMb2mi3xA/Z90FEU3Xj
uQrcGrPom8pyR5E+2+9LpynAldtSRq8Zcv5RDP9JX5UzC46Wz96g6N+mgtkn2HEf65hkGMeE4lHl
7QkSgTEPQU95gFeFdkSbRIzkbBuFoYeLSRg+C2NVZafssUKr+hmVdhlxpaBI8H/Pm8bhBdMuTDXe
baF4PjmAlt+jvXOW//65RpWxZIA7UMjfPM0qvzyqNa1pxutYSAlv2o1PcmRbP4FWJgREZrqHDODh
tH6WmdjzAX/aekH+OByWGjNbusM18D6S4LlsGX3TIzolLYTrISa2x6rD/dhMH42XZ3f4Euhx3p81
JBGaLYR0T6RDiPaxX6lS3M5S/iCG33e7TN4pN6sgdSsnC1dGZG+R0hxlKTJ8/uV4NNtzkPA/n3Zb
V/Ygx3XbsyC5jh+IHQvpMLdvbbZi3eiwvHwY5FHbhbBG5/UA8B1WTNIozV+Inb6mH6Ql6upBbU7n
1BfBMCH3b7kgLpqj8FycR6TbdsifLKegykv4rvvIUfrFos4NRkDaZigtCaiIZnVXVpTO1pWb4zif
EgNlCkNstuHrqcoEPD3crhgsmeH6Xf/rz8L/q1j9Kgqpq9qPUwUmttjr3ADtq4sTp8OgyDp2JaY4
6vYD3iIlvsrZsntzpWMm6c9TPsd5cTVpBnUWd7aB7v0eMN8BEbrJcwZPQef53ogY0XqPYaEL+gko
csex+bKwfWUBCIa0CQFsVSMTJe9XfCiItiSDI5COuXus8rISVFLgwl9d8kiYz0wW4Uc5/jGhwGVX
zhQTdRp0cN9HA57fWmind5vjXwI0qe9yRK78v1upOq1Vmms4KMz/teObjCkPbX2B9HaUQiRhVt33
tNliZfjsVNVTY/oHA5nCz++NA1vN4U0qKQhI2MagqKVuWvCmdyqLP+lf8FTnYwrGXYeg4MOZ0T0T
WzhUhv2C/dNmk8N6/bBUkJuH+WXhb1pveUkLBM3M3YQIYKbjMZTNooiG8dvzTIWbZRipW0rfltGg
rxX98Xl4nw43GXLStEFK8zFBjSoYFqVRMrxgyT+1VKGR8kEYIam3L1ZeP2qWvw7+Yv6+8rFZzKeZ
fVjENVwZ+10eIBH9pHtOZtC8NMv9St1efR33q84L3UZ9YoN+brKClkspTGiw7xM6WMZxur4Xj5K7
3Ct95Si7wTDo7hrfsHA7EZhyCAu3CDJg30Yc8iHhD6oCXL5Jbn4cgi0JAiiIUmXu0lXra4o1OrJG
OEmhCcpHIaRtlsDuyhat8zQI33wGe7LmOThpLb65qT3WWK5DJVxnJb+BNALWwz0bNckMVcWjPjvZ
wbWRKCo3RJNQXFiYWGpDlujc/LoTckBnG42+9RtV5FteQdb3k2KWxs+EyDzmWuwJzt9tmff0eZZC
gktiPz3lhmWywZtI/GZY4E7D6zOo8f/Gou79Sll1LmKjrJoYerB7+BHDEkWr6bl+uR6LvuCO1NMh
8G/+IcsgDLbpZB5T0XfebVnp9EkfVSklT21oxBixgi3KSFOi9eWAJp3zXrTY4RlxpBXcMTr3gvlF
chOj9VsyNQAX9jp8eIZrx8UAZf0uBe5I9WVQ0cOGJDdwumtgdvmAwYyiHwzyGNZ0lUMkzKNMQtXA
2Gf0xVP0mkRcezCmiqoFTGu35veszVCnM+LYQe9Vf18LaD4Cv2ztI1+RjTTn996RNBHkUR0n1ZVR
/JOkPTQGZ2I7wRc+UDlZlZgbyPSSfBJJjoDBUuNGacDYSB5RMhrmKwpu4ej7ESSqnx9xiLQRCJ8k
mhlxgHN0L4RyNYLHfuQNU12gepUGGjy8CgrLxeV3SRDIRuWqMADgfDgLrypwBqPorM2sMs9ptX68
ktZFXcwxJdcqo7diINqZGmGrlEIfuh4cTGp2j0BMfMgzbeYUpfaMOC90U66LKoub+dp7aaBdyyzX
OSl858zl6Lw6wD+bMtiqGboc18KwIF7NyesiOte1SF1CjCbIawvMNlAO7ORmQ5RZyOUKgnkOiTBO
3vgakwZXogeXnYrZXjwAKHlPuWAmiiXRs1sBu+slXY6MDMQv5sp6AAd4wj5DD47Ekvqa49Im77Pl
NnCFOod0mtE0+999pgisGX3rlFq1CqsapTgnX4XvsCrYQmxZsdAdIbjiQxIWZZGwy6zAFPi/YY5+
l9MTHXZBO8G1+iJtEENsF/RXb2fdkDj/p/VhmljDFL5DsGk7Iuk+X8OrazniOoDPqXtFaPPSb8d7
o5CwXbtQMmuthC+kjoomZmrJ7SmFneiw9p39ckPoZA2RqgYsWYTMD0wcwAsTHe8T32VGjAxHXb4w
vTIAVNH5wpxDKNOAodjFMSwz3qBcghDJwctosIPna1U3oU6paurBSDH1fPESGHShTsuCDPkNt/3A
ymgFnsOCYBzu6zuo/jECemOIMVLykEINTED/91fxnmmgmX0J0flYvVtq4MNZ7qWX/Wo5ssrMIMkz
+US0P2+t56X9yc9EsClGzRzNJdSAzFM6c2jZIz+p/VjrgKuyT0lhQPWEw9G2WUpB4xTtPhTsjQ6v
mG8o48RabcM9zOjLqYSQR87B9BHH2pD9pf5QtXTDjkGO/b6++aycn4oNCN+v+vrgGJAEHC2N13cW
RRh+i/1eIU5DUwBhFf5WegUCuhV5e1aNoLzmgAGOTf1evg5y7IJfTgg0FsnHXgMwBEYgCtiAEjLe
0+Fs1Yd0yMMl4q3DKH7wVIpZQBeYYVM+ENr8w9U8jS8N6q0JPGSbCNA3GQaqtZvsL4+RiJrXe3xr
vUIoMnxkHHR+ix3y/23R8hvVvhnvOnx/0YIB0fBy/ema0AnH+iBSjFaYLM7vuJvyCr4Q769jzT5q
u7RGBNQo8mXXoFmEe/suMcTSbeSuK/hwYB12bAyIDoaLToVOhHryyR514+pQCMz5KgS66TV9D3oi
a/3e6C0Og1t4KWg6it+TGLGw8RGJPh0MXoqR7y01no2Rpjs7MzlLH3E3IYZambc9YpdbtDCasv8W
Q5wKK2d9xr7MAU9XOTwscE4Xv9d6cr/bfirH7Lvjg2LWz6KWEu/UAn0YQZ+V/J4VsTn/bVrk/eaX
PZpSsFSesf7JBcYVGbKbmSTCH9iYA3dW//LvyPXuTz5V3686tABQqe521AR3OcVGr/2VHkbt1upz
PvROv6o6kNCj7NZTUGGkn4ZIjnqqhPuDPqHlVtHGN3t0V02WlcB9gqiVB7Z2sGteiBHKp/yEXja4
WbAWTDyJ7DqA36BuJwDo3vAQFDA8/dAvepjqYD5r5VqbJqudRyjsHuOLEKbdtJGZm5zWvGYYoNw0
ARqR4aiIMMSp6nIJUdiKc0lWZuie+ubOIBGZoX6OjWbm6NGTODFAD61hWGFgoR9yL7yhLuMtcrGg
1TKst12FTuVTDpT519TrwCAavJu5jLB6vVooDxUWfZRhgJOub7NYxx2A4aj95j5s8TuFqqdLPP0T
H41qe26XL2EUnRsQDXFX/JkHH/mNpXkNxNqJz/c7h08UTGn0tsEMypIkGYBirhZWkRC6YBrKAjzJ
NkVXRmNFKCPFwh7DsIYwq0hUjS6fd5KB4Sh0Go2a7t9nBhMVMr5R9QHyQr/CGMKLzvgpaxXTpHR0
mTkHjJNAeWzNVdYzTWG3sLqhC/9dFOfU6F3FLuN3WlsEkpyv1vPQ9iGl3MND2k5O3dPIxobPRmf3
o0T1oRw3gEQ1Kj8777jZO9I8Uny3h5KOv7pbKlOWeCjWb6MJ6N4Ct0TDBq++Skyv6YJipDIhJKqa
pL9IgvVUPM9ZtveUpCFTSnLh9WPRuJOTkQoYQkSpyPQuk0z06SOUgBU0Oasif2RC0ZOhOUlalUQ8
iWlh08Dv79eNGZIHJ2wstW67cX6d2mOR1u8UerxZXwuOWv9t/tKoUYlGruZ3JQ1LwWVlk4y2K7/E
cXY9I9YCQPJrMV7+Us2RifXM900SRft/vmFecRAQ2L1Fw9cy3hd7YRBcUpf7fL5s3i0a11xQQxXB
fKiiV+Dg9Xj3a7HX/u0bcnQ2VDgemdvOJMw2cNl/Q5S6zTYjGpvaHwFCd/46YWACiRCG/5cKoN/N
ueBzxbkXfVAkf9VJNTy85ep1a+NzjfuaU58ahtvTO9miRK2ZbucCsOeak61+6CIbB2es45bLzRml
6xUZSEsRZDN3t+uvmw/ujPADTmMzltXFpRqu1MmSaudaOK2aDXAZJj4/t1SdaNwAi4rMr64MWCvM
8GSpZVXHAaQ9MRoomQALFHzCNXBftQALac4Vm154Rr9JdfpO+C2zRAS2zrv0jBukrxc+kjOwKyJ7
oAKfYroPTvkgcIknimdNFqohPzHvcSroA3qsC5aJ7jnQEYtqbko+0p+U6cC1i/x7G72SPOr2cWep
jMkU1vNJv7a30OSBx4zak5x6FN78jTeGb4CUaxVMBVHzpYdqllvYP+7PDZeZ8IJcJb9VHzWWL+Vy
SvQBtEM4uwrUSG6Bo8Ecj3HBEktuN33NYSeSPXzzuMySZdAALD6Es2xXigIVqPCQceUDCVOe3BlK
WHF5B9WHHOL1SmhGO2VBaGYunZCbeQdtI5p0jnTVH8yXQHq4WzNk/v+igL4NWTOOs4Mp/prj+wkE
BCttwh96l3EqP2y27GcHnn6z4FYKMueLuhDDh4vSVAReMFkyObjkr958tFwKukAg05mM3Pgh/LmX
3PzsF4PQXOQizNvIyNLkHZ3B6iWi8rtPs4KQKEu5ZOsbQC+9
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "P-2019.03G-Beta4"
// Program "Synplify Pro", Mapper "mapgw, Build 1429R"
// Sun Nov 17 13:25:13 2019
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\e:\gowin_projects\myproj\myproj_blue2\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\e:\gowin_projects\myproj\myproj_blue2\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\e:\gowin_projects\myproj\myproj_blue2\temp\gao\ao_0\gw_ao_expression.v "
// file 8 "\e:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_crc32.v "
// file 9 "\e:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_define.v "
// file 10 "\e:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_match.v "
// file 11 "\e:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_mem_ctrl.v "
// file 12 "\e:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_top.v "
// file 13 "\e:\gowin\gowin_v1.9.2beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DI4rXVSqQQakdxUiFbNMpUcFqLtxiH/v9VC2fotO6RT5oJx4ujfd+d8ntglwi9SznfUhuCDdANfH
XYMgV7tqilOQ2ZawjyjFzCrZ5SPXrGgsruT0nRljnPbi6qkiFtugOcQTRLawx9T7//cBM+KloXTA
NW5UEesUVY6XIevfIUZGJ1ure5Ny3juAG8DwrfgVKoVsVbpFHGqkn14/CuCrPfgd3cNIeMnz2tdU
fIIQcJuw7/y7oxsPIHnSNjduB2VlABUbTul3/U+MLlIz6QrQXnGGd0gsk0VzmjNw5t92AUKNXFJQ
KgZfLCLpjgQ/ZbGsMSNTxIFdLQdlxHMJmC0vaQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
BJq830S/kOcQBA2JJ2q4S6I8jB9jjQ+2w4M1vD4Tqw23sKPDOhifxjr0/o3W8kskkjrPH5ExmJnx
4+Ax8NsC3/y94RfnMYtaR48dVDd/uZPC+H97z8xQbMlRtAPIPBxmvbm2XF9esKwvNQk33qXslMT6
Af5S+VRtkbzP466p8XNJQwyztsU9oaM7FXV1jV3HosbJuRzcKVPEOmo4Dn/DOSxaP8rd5LPjoLqS
+itgiiOB0/sBM3oF4lMqNh90Lt7h7dN75Xc5z0AOiCtIi7ReGbnoPIxpLrTX3YY2f7/TaNJjwe2m
A2muDv33kmPJYj0Qn1mVE7WUxAUWY5au4KLJvA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7376)
`pragma protect data_block
3l2m8UONmp/7H9fdVZbpxpmXcLOYUQ8E9OKnRpvBGbifTTNhr6GEkq1w2IkyLRm6yOYZRirjYlSH
8jOV7Wk6V705VR/MIi9T85aXx4xP22/JcuLNq+Z+KxLcZb0lz75Pr6xxFavJ5h87IMuWbOWvueJz
fBVyWZ/ut2kxIiV/KSLIGPc6qxtscLPNg95WBIhrUN/kuNL2vlWdH1zOqrpPeGZBwi0mspOT1nhl
4hjInY0jPbmL5qPUmHpOp9/9bquf8Um4HqCN0CEArjifPkXhA9yP1emBrCPZarXQUKHvB/glHOzs
SlKgEwHLQwBQso7LHlVOu5SSlrdciJMeCCU1jqUJI0XcIi2j3yLDPRWnCo3XO94tLGEgCf270kjW
WgTDAMGFeO5qEoMvMnXzc9k6o06X4W8uixawlyxG43+ZBKbDN5558IsANrQpBzwpMvph93iQLh6J
yEZvF/vUDNaBpNuHMZjbyhVBIX/XUKaos+YN/tyfjR3Un6Fuaizwu2vX95edJwuS1BeTMMrVovhu
lQlTCAsm96yU3/yKXQuHDXKP1rJ4ogMafBHOE/oj8nVqo4566oVjxnVNHSuHBXHkk+Xk+YOWrAMi
FYHwnWWwSscu+rOfpBWCGfNndmi2QIWyLpYkVxXpWPSi17aU4LtkREVCAusH4IUqgepUMHK/uS+l
3VubiVwx1BgmFNXDekVkGX3SfLDV8cmvmEEwEHyWjXyyIjs5Y7QTgJgfk0oaXxn9+i/m+LDRs8r7
2c7f201xo3PWZKNot2MVx0OVF7Q9s0PgYz+qPlSlzPXGUvmzroTnNLhkTbv5amkMVYJE8sm5Gr3q
Jo+iPSOEpoZVccWmE9t7GyMmjRzwlnyWgJ2uOXiYko5NR3ks+gJ3ZmQ7WIbxwWIHzb/czY96kTkC
sZ21muSILD7lK12SwHA0xaC2IGIE2WZq/jhVjky4PkNJKXVAM7loFa8ZBfrt56kWU2mvfqiKOsrC
KoYfnX4eftfTkpQDw/nkJA4ZrBeQOk3tYqrMMlJGKcaIJXHQDUNhZ0nDF9NAwgfWYolo2NK1Tpww
o+N41EPUGBAKdGwG0nUUM2aW/lNoNVZ8dIjpCrgpBdJfuvk25+0nvPqdyOKynJNBEWxdwksUdj/T
9hALxYSWey0hciJkw7GBrTcYFcF0Rqr5C4wFYThOmW28hzuIvnqiLZ9vUbW2lnYh7y3B8Kus2cCd
TR7lhXCFH9ypH5IBL5fteA1/LVyiaGbpkzYZ++/pifMWVS2+IlmIGjXh3v4RDuoAebqn3UdmNnd0
kPhl3FxNE7/am8u4jUUo00gB7JKRfQsk0A0x1iRACwxRZ9V8Q2HYpBmsbGL2m9/EQM57ISwztXik
b4fMvXNqVF2ja1kAmV+sng3E3BBNIQu57d0+aDr+c1sYCkTQ82IwEdkfBJsSMf6hX40CknkPXqmw
FjcFjrrtZO4RYzDu+5b/syGdZo5RpJkVeujET+z/ADW6zkr7YhjQ0YSKm/5PqhBc/N8QAVbsgUpz
JojpDf0Cck5weSL62l8L/VwZ2hyqn9Sjl+FlOJn5Pk6aSdX1ujHYJxtB6Th/hv443KHcVVL1xdoI
MHzHLd4S21SiwvxL0WoD0nEe3VZQeFfYWEWgY/LZLCAwFWXhYF7d31FVPgBFUukEXkZtQ0Ml5TuQ
4rs1lJkHx5BEEdnckjq53F1Y0C6i04gMdx0QaBxMxQiUzYtT6vsX1VczmON6T+LMpjvEL1ITWFKZ
LOjMoUUGNRlQ3znBqSx5ZE4DCztd1sE0VuuuRUiFbVuAsdfLkLDaWYwSn3Y6V54xWnY+yIPzuwVU
35a/ucSDscb6Q1BFIKTqCI0gPL/l167E3FMOuq+cTAEMpkdf3bF7pkBBjytDmrSZpKSzxw4zHzL4
AsFdOC+zWKmvEIS5Ipt4ktMGyRo9ZKxsul1ptkrJAmWgjjbEB/2Z9m/Q3dcPoxg7neJ2zZoFmIpZ
sWE4ztTiKyUojBe829sU1PILR6CJ7XQOGcyQCndRht6zE/isGeK+a2xzISvQ4WCPGOOKV7wxBEZz
Q3zh/65vSvQbRtKgcdwjcy0ZyGV1daaT3lNGblRCunB3EnpvEtM+6CD3O2hmSZf+zSV7Z8NUJpBk
pzcPuU/9h+9b9hcLJ9h2XxGOGx93KL5V82UHKKr4UW2VZQ70h7+mNDQux0CMV/2XaN6GhBK/JcwH
PfI1ULNSD9J3DE7gZRvrHVOl7DvCINpkWDVS1vwH9I7dsOmA8Gsju4QbDTFsOlNK0IY8bfZuHTsY
7kd7wUUlLtUSiyBnyq+TAtDwlLZN8Qy+jLQ+D0uo/5ZVDOh2B9mGeySmyKnyCdXNxN3SFYWxnITn
Fkp3SommCMeZbbbpiACfQ+V4ejMZOBoGt6z0eQhGC+2QL+SQWR987HHXI455bi9i4lLDaX5li/zg
+SkroUpaWZh+2HQeWLZCBNhDyZWPMuFaPdPKb2wAbXmE2te1Z5Z7Y13oKXnDa9cd90rKRqoFlUEh
u2tSaBsRwNsvl2yxP8Ai38pPpShDNEGmGUvhDbj17qE7ocOgFYwNMwKC6b/8nh/B/bZeYFISDNQi
vuO1m8vTt4bkOOEU6jWaw0HigsSNLC0DsMI9V6b6aRB7kN0f6kLIdFfN3rz+NXoCaP7G1SavGoVE
UEPratGEAFoPSd+7aEbdgrLqBELF4R/8b16snElxbYEM9I+k+ry8t7KqJrx8C3VUHW008RHWVz1g
6+UL/D9fduNEWhW1Tfab05WOYYG/d/z0S/6c+K0IBN1rUFSb0oPFeCroLdZJAeX/OH14997cBIEP
vF2bfDOMzGhUg4qhZ+gg6WEAQgSSzYNuThaCmixWByFrvP086IwhWF8Kc8YF9VBIrG/FJANinv/g
r+/+tGjwiTK35EVH1vcuAqGZiiY26vcBW/NfIgtWF9MSZualVKwmYYAMiZD178rUTeoCOSnDb0jv
7Vok7MdNBOFgNXDGS+DpytMpR1z52YjxibcNdQllnE1umOoQDUEFfa0yv/Ppa76oBo6yATLqlNSu
DVo2RlYkFfhW22PdxmxzDX2K0JKfJvSj79QDtO7VWNYACLIbG8zu0QvyuFLMAZPsjN4DkrjWm861
bUE1tDLoKVfAyqbpSEHw/eAmaOrFyvk1BKI5MUpQYI7M3Uw9KcTipCYbJAVtWKugYPHpdiH7uR6M
G8jX8UROcRf7MNF2x5MSo9Yng0MYT/UhDFt6NsZvKgPpZjTA3ZmPBLW+awa65tdZU2ya4Jro4WQf
+UBWOhxyDuTmD4MRxSImvXye73uvnknQAfr0FETl+IB60pbAgakK/zLRBehP5HhaojiNZ1fcDSbo
hnEIzwsN7pHfclaenYr87vfgFe0+sjIcuUzxmBHW9RX5l17EaSC5exR9UB40tnYrI5+/ftaUaAUM
+Uevmf9K5HzHxQlphx+7fZrSicwDSFsUB4AoBZNzv8fpt24zuuQ+wqH5Z/7qokYlyuibPfK6SWBU
+TuNRiVTmwRoPDMM3UqTSaKYq6BhjXGspsSzDp4LV+wzCXLzhKKxIIoLAM+d4nS2kkTURW96EamT
IR8qPmhQkXKQsl35f6AeKQxLT6x7OmRYy7DgQ0UKnMvA8JzTXlhsbUHswvwfio3uN4/DWf+I5RyV
57hVK7cJGspwzr1Un449d1iAQPiZaELMjZQ1fAV7L9Ptkb+r0KrC87yRYmpgUD8moZJC2aEh8ONa
M2YPKFcU6mjfK9GM1fSCTFZl4LUpdA9dvTeEPED0bRAtUD2H0gNqywlZDOLVuNGDVcq+oF3t1egX
MkteDFml+7rbCKbEyHBIoIWI9hQoJcJkuyZrJyfnf64Nk+I05C4u3Bt27IgFZv0IFMkn365uP6CV
4uxJkU1samkh0jPQ+cYvpdtAAKVnA7Sh4shker5NDEVTK1rmP/l1pC5yFmNUBQHzzHUiKYDIGp0b
qT9dZdkjZPPJKFHMK6LRuV6Vh/eND3+ahbRgL47f+ieG/vjnSfUaqiefLEw6JKSW7sfA8Q3MDcZt
/XHPpwuLhIfZPLId2wBcWp9PvcqhZzUA8AKGj04V5+/wuOkbOCuqoeMPxV6uiM961Mh7yy+ieVVm
Csz2ZV4bRPagZUPWoSo6PpmywXoFplahN5ZJkLxYFMxF4+LXxHOkNXJuf5JI123j0h0lA598UxLh
eZSIPmv8tQMuxEsxfzIHPqH5qcUg79EL9yupwnsZvutl823gEI8m2B/wU/ibQPHiI/SkeL7mWuPr
u2aTVhiKXvcfDqhrPPis/Dp7fW8N2A3GdPj4XgK6xlBgYC85ppmQCp87SlUO2TVCi3F1mB1hQ6aY
B/mXDSDYQnD4ovUdSjZ6uhBOBrbF/yGorjo6uTiY4vuJpsiGe3Q6dnO53GqWfGgo2dLyaMK3uIdB
ECrqdM8+Vr1gc85gRZsLKy8PJ5oSUoMyZDeTBJHOWHxPfvEi7gcWs1N8mjdV3RdERGGXEbQ+K7q+
ufAwCMFEm+BufS2uSI2dEXGGvw6aJCjKq2iY44bh+SxRfkpLdbrl3lbqImG9O0WxaIUt6j12o8Xk
HNI3MS0PYOitbt0na4ipfh3vwjB3IW7BFMkvWqA52eY2YvESL9lH26PzjmDVZctcxghhCw5bD5mB
dn2d7SfQauDfrRKAJaiviK9QVX+hL5Dzq5cX1lVa3rhMT2RqMnQorlKZzUZz+UxZiMIRDHFPavTV
m0/2fVxOXoEha1Akj5Dvh2j431UYO1FWnPJ5DAFHp+8IQFLQtjtDuffqoxAAXF+0SD6d+m9RFGFs
VtONvPWncHSyMY62mD/sufT3N45p2NKFqa+O6YNQJgEbiCnjcMTa4l4Pk7T85+89JO1ppDaMY7Po
9VZkq83x68gEMsDhJCi1+//F2P7yBvV915yZUAm4w2HcXW12F04Y4JydoIaaKaLrBx9q7hYpZ7oK
ZugqPAYG6yY4Kl8KBeeRPZOnYmE11RZplbg9y6jx93iceaUSWm2PbrKOAglPJZ8LywgFkUA1A5eV
6wDNRcLfnVezvY6JsOEKAi0C14pzmXBQHZTonqa26cZAxE4XT3YyIxH5XS656DlnKqS2mQakVhTc
ukU+FdhWLauhkr1n/ZhRFRdO7XHKZAk0odwQTCsarlrIkEi+SDyEWJv6VTT4DuyGcsNza+VwIVoj
wBGGTdlJaHLzN859Fe8Ct4n/UnMwGaq+xY/kYMwnS1/sN2QvkGgHXy09nONMVGfEkAXZrWr5xY6W
tx8J78I0Mq05wQYOhmAh3r52If8Oic+AN0JWBCuH/77PWCW7lv6UYTXAm5xuxeb5m2CZ4LAgQFMb
8FuJOzYUM//pZYdoya9d7LX6SCKkh3l/7m59xvTqremyILr2xi+uebmPLlhVHy6lADlD1Ke00RXO
8JEbEGJyFaszdHztBxJQS3EqRu9uFJzZ5wm9MQOdVWEfba2D3r/Z0dkpkjTAu2qA4QgZbEj7jnZg
gVaEKcW7pCPu1ZTD7WgKoaPZklrR5E9h26aZqbSu6HbCe1fZHJZejgmsalJEnFfAHlWBn7ZbJPaf
sNMEKSTVdVHeAX3Vh3E3qnQRHL8zJWfeC49WEPOkFnxweQtukZnnaEB8nSLsoBmV5F1K1vi2sc1w
kVdyDwamEaTr5M7HfiXIWj8o/s4ZgVWCDBHKQagv7EXaDI3v8w4py1eQoA8zeLxsH3b4JVMGft8E
sKYLaDpGDbDeCgLleaEAVH0u/1PMfTCqAoSPlVlQDOBcdlZtKv/+5fDMDZ1vV1MZrR9CGfDNrojr
4DqO57XtKbx5Brt9UwzEfdItmKpsjyJvUBKflR3d3O2H7WOqJCV3p2oy/yZRep/G4AnOCliRlYZ0
5s4o5kJPIXckDICECXYbhGpuhF+mLgFbjP+JLtoZTVO7x0ehzrks54xwLq32xNSzNcpJ3gsoY2jv
3ezYf+xc1T74fLBdBMwH/iGTxhztJTRijMtmkJKts+MXEPmxJmdaVsUaATT3xRl6mBlXyyTxKaYe
B5U60/7PWMhbdZXrH66scM6j0FatbG2ZP20xrQXOSgJjaWDgCClqG5BMRMGIS28BgaV4qzW2ds1L
KkHOIGtLSZaWHX+fSmxQj9oeg6qIwcv57M/ndXNWDXXGK1SPDCF6/bYJP8yInxVHUdOlGDyPXHqE
y6jawig5f3zwxxj4JbeO0LNZxFhkvqj3S6CvGeBxqJPqdJwPbNfZ+cvwvcSMspg10xutU0ff7ZS8
8bwFf002/Ia2WXAh1ytfU1Ss0rlDB7bb7DGC97WDn5B1jm/WXUqusXog8Qayi9vJq9lVZZpGQGN+
pA/rpTWF1wNbl0iat8F/C/MkWUyfNmwLmWdF94xHLasQjL8rF40Y/WzI8XG2N1vVhabaVPOxsQpn
U4eJyfjmHv1XilXGGCIVjf/Du26cPx4TEggbDFH0qaR4hXgKPRWs7Wg+yxxsxu/a8qIz+enp3XJv
pAH94ZdEePPRYoO6dsHL04NNRtE4p3ijXpq9V5cgGKLvSlrioZKtfTF+kG+c44Hp6X01QGB8jeMa
5hXLf8EKPa/P6Lm4bSu4i0dEXWWDpV87nD6EYzMoWYkO9fxvmTVcpEBozRsLjDDLu0zEsCECdUzl
ir2MrSyDONEal/86jelvIJxDWsWxdyvpJPi0OLFoTtx195ubFJXbBF/nqA80qRbPfzwIpmq5TFZu
mx8uspbPlWLNK7CVLX8kWqBnYemrJgDjK8hXKAEjnTskZ/BwTdXho3IRDY0b8aJJpZJWmgcSSEKP
y2v2YGxI41+0PmEmr4QSFXC71ZpVl3wAFMfvW9VQb1YWEOFY8mYIdyiwgy9UbCSUqiwQJLBvMdHz
x4mnYFX4WKfrUAPsJI5hZU4ewmNtOQL3jVNf39E2XCGC3BD+VIP3lg/b+0obeCTcKgvwQgSxKce7
ZJ/B9KrS7va0E37/B+jKZLinUQhtNUXCMUURiSJVqR2XjWZsPA40VYxGTanweVkYGfh5kMrOW8h7
RS5AWqLNWcC+7piqPUvIwb3kAPtMcMZjB3rr+MBU+jLjrusieIDatljsUxuMZ+XvIyht6CFcE1bg
Y+82wjkHfDuDgdwo+KxQVf0SGztbx+8VbcXZV8ba/pZjaJxYiAUNcdfiugMg2tModRG6zSjm2bm2
9D92uhRBIBz//VsEt2LmzssLG5ydBfaOW/MTJ8Av9Mq7ZjajA0As/ogAjvWTr2xe4EeYY6as4yH9
opllq6Annc0Y52liJsf0IvCRM6eNkRQwOSMd6LGvvKT1ZJs6bTbv+T851FFwMd45Do0KZzw6VuHn
umi+aStJocqb3SQnMzJL/hYe58pCW2RtCZIxhjoEqWnMpVEkam8BMwGdZ7R7rSLvPzbf4wandXhu
gtA7hi6h83ogRr+FzOMCSZu6fgsVFW1LGu626ODUrhxVoRjkpiQa4H3Cp6FsJeFFquTxKOVprcRI
JKeGExVijb0nmIeYudYHYkTU9cCRZ7JxnY9Z1BBm3KS2i412JJWg4/ViPv+c/wPRA4e7y+YWTVun
7+ZH73PUph+Zv8ux0ou2ivumphTs6FGrso6vecRvavjIs9q0DG8hKA94P2+rke1SaDH1t5YIXMIZ
G5XSWYMOkGeRCIzHOljOVyCcx+ZIpEJXDEtrQ3DFm7Pcv7TWks4KwoGzcAnzArGxaP5XiFWiyds2
7kASGRfjzkrKq9fdE+broUxUkP6xdvRhF5DWS+q7itBhS1zN/ShADIFOHrWIPG367wLIShnX5Mk/
9lD4878Y345AFYYrfA+h9htoSqKO7kbxUtYdOZkzuRHUJksjWhiZ91wOvFZSFu5GliQ1bd15OX1a
euXhKV2ptwFufayqCG4taaeydmwaaj+ABcJE8JYJ+ShdzIBlrJcBYSRGZPuSMa+J2XBPq5c8hP1d
5Pr/g4t6R5x967taC82LbgZuwKnDhvtZebjRf/42RI8rTV7SBtP8UGqICCkvMxVzlbzZac2Kn76f
AxppbdmVRhEcMA3NEGqz5KM9jAdAxJXukTXtlHLaYCzw7q3VZmwfSMjwnYiiqaggEMigchS/gtYT
bDvyvfAUX67cVlFiLDHarA/wlawCnXd1GUBoKLalOrXAx4hO3CnEd4EyoWk6u/W06cwUAwo2Xm/6
c858119IBlqssYSmPNuFm4RJP+5epBu8SY3DrWnzS1sbNLfEDUDtNT9pkrPCIJUnWDJtXE/WNFd7
kzkb6RfO3CHF+33BtBKM4LM6u3oKCh43uGEI5qZOC+UXyDfB0obR6DPWxAAzSUP3o/4b6LzBu/db
JNTuC4QNQekbz6FMrz3sINTJh/Ea3lKXn+BO9ibr3ji1cnRJVqsyJl5LxIxWHr5uEpIcCJs+J2G0
UtsLIc18VyOTAPGYs2d97Ufv2Z4Z9l+I1Ze1WJnIx5hkorGO2xpmMjBUY/+3cYBmHRfNdAbge12G
sHwHGT9FOexw1qmBu2Ms796aiTLmyFvxLOqnKyw/yJhSRv0VoqflrIl89U7/b+PDHCFgKpH+K/yr
aRCumf9uALg7+fBxIFJibRX6yD+K+4hcoHqrlbFPIMY863tHTnqncmM3d8dNxgmuK5uOev9cplYO
AWboDb18WpkacdgPbUbZYPMM+0qJIZ04+IYyzsy08GL/Y4yslz47XXW+QTUjdohdOgmxPLwbFHjO
/y1LeLxpLzI6g412m7exPk4/9SHfPZqBWUVh1TI/GI9crwEbMpxiO3dcEN1BxbdONihT3MFKtDr0
DW2+/JX5LYDguoyzkChCcUsQ2gcw9+oGLO+Fzh6pWIl3/Jspqbm0CcivsGdPFK40G2lElL/VPJ80
y0zLpigkvb8MXvFIBkZeLSLLNHm5IW1delrCncXJFS4xNdWR4XWgxplrqTTkF/4GVBOlO+9p3p0W
oW86iVl4Pf0tFvIFICJdz2BLysFBCrJA3HWuzmNSVJ8NqrVJRzGaXDt7VABxpux8oQU7PtYWvwUA
LGu4gB3JpYzKyaOAUH/wrQ0zMHYVOLVC1cxzCL21wJJllkoYZLW5qf/9z8teRAmHgfr0MPLyciGi
jMOYrhrYEuHOqqvwwzdgZFl4uDSpulnXrSCvDJGZG6vgQHCZx90+fQVLG0TREYQbpAinx0oLp8zA
i9W7KJGQMJwUeN4CP1w16nEskOwQoDkjxGpJgXWuvWDqIrPqDMj/ZmY1D1+PgvJTNdVdoZ8gCit+
HiJAWrMp6Q82T35WFjyPyoQWLL6c/MnabLDtaHsz5UHeVwUpwd1Wd1hjaPyRDHThocalhWrOn/k/
cJChlG0V+RnJ8Wfg0rfBb4oqrfXrQTnMN6PF3dj5GJo6xdWIDVBr2WbDKXcdq8PxkDu6zi4+irZG
oL/6AneJf+CHrbO7KxlTSGePQiwl27OcJnoTgRWq06jks1kxij0VylkKxx+Ejea9JWEekx0hO2qU
g/aagBS7nPMIqnun73/yOU2K7eC+o9g9ge+xsh2rGgwG/3EfdsOanbfXOWv15JpS258ugBuszKh0
SsZ9NVizbuR4Ls7AZpr2/G8HbkU8krBot88FoIRfYnE+INHKIoPv/joKsPeMt5NqWYdr0ZmMhLYs
rfKgu0uEq6M4cNXKast7ebq07J149NGXNyujGF/7LllUXWNZdlZz7zJFeM4OYqNBHiKLBh9Zkdev
l0+Uqh+jNQfH+pTJqn5MKJPpl8rZEVutpjfybU5EWBjirB6lg5LScidmGBeApGHpLKhrvPubG65v
FcIG1w4WRjJh3VdEUdGE4vQvOTFoP0OnDiJCQz+dptfkxL93t3xFDdne6a1gC7UXdUA7ACPDghf7
pVRI7OUFRBiu8bJtifNh94EwjXuDQFg=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ga7z3iGMhGhga7TzPGleypVOHJn9S7KEP16RJ6j/y4QGRddc7/SJdXJ2zPvm8FTCqWlJhu6/s34X
gPP3kw7dN1YdiZ3wZ0Vzt8uhC/B62KTkMGylsJT3Hm/4AVsby+VuOus10FHgOgp78G6FqJDW2hD4
FEF7AvpJ8kF9S1ZR/yBaB9R5/vEzgMTG6H0b1hzTpBGPyaW1S33KG60mDs4uY1wSc9WkIOuDsX13
gE5v3E3AdV0s35W8mk90srPFan8A4v9WhQvKv0pRdTPwajKYNoHYw9l0a0ijfdCCo0SwbSJr+KOr
7KJQNnQdeGn2Y8dg3BGFPO1H0k02bZuSqUQ8rQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
dBwrqXpaPIvc4b2fzIcAYNKycDBKm/hw0N9OirP+O5J0w47WHpIJLrz+YZdtlXZ+W2OT1CCdKga8
l9q6LpHNXfMJe0tSBaUQJS9kx12QCBYd7pz6Zz4XteULmwejqAW/r/1SNtjKdsFfgoOhPbvsYv0n
RR9WE79+rnvNSo03sWloLz3If8EsTQUj+4AuHA6W5eeLCFFrjEJDELred9ftNf+GjbKQ4DD9VT1l
GYpqKI157tMW7VzaYctB1tIYsZm6N1scQY5/pen6aJE9XG/GVJc/lUhiKfjKkAB4R0V1b6xO6o/L
Z0CvpttfY2ekIVc0VuCKq5gMTfn8BkW7RjZNRA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=9072)
`pragma protect data_block
3MLlIGXYAu+SNVZUrN9axPWxB76fSavWP25CyQigoZQ3T579rH2tX4mOroKAFnY6MCrE4zy5SoFT
o9pFhWobhy1JNncmCcy/a0fRL9ZlIyjwjHAt323ZL0R5G1zw5cvTmFWPoZX0yo775l85Oj07XBYY
i+0FcCRCKdgsQGwhMUnpc6ET4ttBmjQUuxB6g1Afy5ISJRNYs77D5E8aOFrmzUzDFsE9BGcX8wUT
bT4zFmjkBZBQ+KrbdhaUiVbninMVuzKJe0egFOCGcc6CdMPwZP2SxWGkscRsjPCAUdXGIydg5Z31
50m/zUoKITRK4jViYvnHt4f6sELIUTWEwPvxSg4M+j+wpDH8hMQC98bpm495w9Lz7AbFBmLBe5IG
17+sbfU7k0MY2fUrDvsniZvkyXNkbKvNrkm2E9MAmf3uKtqsnMU/tF2um9tYyMuoXrnv+cf1WHME
rcGa/NDEnGr3zL8P+jWgeThli88TgswwgsRldtZSZHdEDO1R1Eb97kPR2KAaazYlo2Q2STr+5F6V
SY1q0ie4TtY/nmeVptSZJNGauW3hhgmAK4fuCh0LfgbkBsnHNuCX8t9sRAwVUkoEOlvg+hIeL3ch
IbMuCTBsi9ym1EZ2NwdIt6YMzhAa6xgt6mL0uQSzppyrK9CSimYyzPbah+kviBaNcZ+XJClYLFwg
Dt034rBFaffea3MI9/T6EckVHZwmBgwvpnfxe5dIdxVZcMCrn14d+8gHoeJtodrk7RCejHv+C9Jn
yRjIaiu6w3mbAeAL4r66PbCB+S92jMdnwdBtSBcwI+pRfl8Y1ZjnMUax1D4+e4G/2vS04zWOHJPK
TAm5M/l7TRLujzCl4M5tq+MN/Sl/TrmT6Z4/ZBXtoFpOHicvprtU+bB6bA/TDiQ+wyauUCUWMDnD
F2sWssLTcUSqWyGH8nZQJkJU1GRznsjpDp4OUZFEoGr1SIfqUXOeUdRWE7kTsTGtuLLkFRULD9ZC
icKwOzgQXLWvy1haIHsyX6SZ+d2z16A+qjc4h9yGuTAjU8NLa0V/nk/gnsMB1qd073hph6QLxLJK
r4sFXdYNYgCk5RaS44kcalofpqStJQULijgevhq0IIAiHku9ZgDSCzWAw3Mr5M2bNizLX2XXA2zw
yD5SKKgh8NLJ62Z1MJq1d/+XEurLezROXf2MzGpmtx5eT+YNTMToyw4wlcI7tOteLNTVwpN45tUQ
B+wyQRROLfJbya1slSCz3CBx0TkfIQfh2iiO78hl2uIlnw7hygM5cDhSSbRATA0xa7ahqhvOPN7M
cHlx2JtFdxdsqSaZD9QoJ639DDyU3Hou+ECwMn0csUSwgAS8rtGVdP0Of14CplgwrGPXstO6akKA
3u+imfQ/w8L/PLKXBmZ4JDbURy7k1H6RKbw37csxd/ZvrS/pSmIkcNCzp/c2DuOoQ7gmrvF/T6P6
o66nwV4BSbtkXVm1Gd6pj8kuzFas4d8qUgIJYtO74n7f/EHBC4KRyKr547xiGiwhk9b9qd0mjPKY
rhYsYy9gXuZh3r68RGneNEq01MvW6g9QFwK1ZOIvZDYOR4QWzSf3jaria7TfeR04B0hTDmN2pnIe
G0GNQyny7szBaDLk+3oC5dKi2x7IBMiFePNumBGpRQwF3BZOBafJAtsThr6J0+IuaIyGTu6q0CRE
pK6/stbZUIyDHLZTtsEiDvCUoqJt1Nwycg1jZabyqczbNym1H0NA+utNZBXESxVE+E0tL5xp64UF
6UUd+qxyLwKovERkzivDR8GuW1zTirEOV5S4VxepjAekJHQRl/DLLebsO05p1WmBlr64t8l3I2Z4
eBoTyoAckywhyY3Hef2UK2jwBO8dnRLD1Fu46o95g5M70RM/CdS1OdLKSF5ccJEDtzouHFkJV1Uj
jF3ui454vNAg2ROOQ3kKuyo5BsEY2EVCu3TpZq4c/q9GQLsRGPOnx3VcTR+6BZb9QBmDwr5qk+/F
Mfy0nKqqzp3OK73AWybRMjmJczTm6ffP4zxEkfUdzR127EO+OljvRItBn8LSuKgqUpIu2NxDCg+f
A8xmKgcdP5Vj8cz+tus1NipaLcnS3rd6rslS/DaabQM/fOpx4ERbftZUSiDhPxRfGlVjhYH1zMEk
pr486KmY6LfVGaqc2pCdgIkuSoohsNiPN8xmmK5O9HjxRm7IYdaUIvotow0YeYsJys+80/gJB5s6
cE/ss5YkBWNMAqtri10qAqP/lHRchjbTFTFInn1auRmyFcN5WTjU9MqXhbmBIpJrVs6hQ8bjrGbe
udyynSp5mkE0eE/e2v5I1wi1YhxlXU/wpSQkq7AW/DgOKirxvaKomORblPuNuqND5ETjQo+jpEPM
80/aOZIyPqN0aWmrTJE0jsjxS1AJ4MOENCzTG523Wq1bgye8XzrN4fo53VpdHD6EPKSh7ZgGV7sq
giQ8mzKHA5CetG2XXI6zrPk7Oe4z8m90oe+OF3HP34C4sTOp/x3Y+GqefIC7NoHPNtvs6PK4n21W
QJDfypWh5VF59VtNEgflzAT2wYDVtih7VEgDNBwrj5ychDhaeRx4+0dTJ9BZTa/Q0qZqOY4erpsq
jvneKxGNPh7zRngog7RWOBuH1Hi9ahuIiY+gEC8RxoTw0q9WCloHfF6cK42Bey41W7Nkg8Ic3W6O
AV81HlRcI218/r7yKU/7urKe8KAq0lmfWI0uIobow6NRr57vlBBhnMIl/DXynMAD0MicHsH1Dhyn
h+XWBoQuDUWkaHIh4zZ/+1qRMEs0NnSiSUJpOxoccGc+tyhoKIypXhHvUevk4IqtTmdXqAG9BJVV
k5OY9fhhlE2OW/ibdkZv1N8TAqzbACTxaJsG4yd9IXNrWQH3memdIJYipNklf5EjC/KvbTm5tyl+
BLxlplNCoR4T5q2klsjPNTl8nKAiMYCZJ29rISm9ghJjvtpxxC7iQxNuwy8DpjfL8Uf4MMBxii/H
GSJtEZy1R7DGqeOvCIAWAjS1+kkxdMrlh0x3ruEo2+mWagYuF7zcRwv3TrcxsdpZpxjAK3KuJQ5d
X94lkof9p94Q9FjBqgLyhEjFTPbeSIdMHrEiuPoqCq/SHstw6UAe/HyD6+3m2O2WR1U2m9uPatvm
sJxRvmVVaHWurvpn1JNRY5/mpZqXlkjzuf/rk4eL7YaveH1F0WX+Ql3Pd0MA4RpPOCPoYJ6ooi3X
oVoBCaBgNLwuE9nJoaTWldtbdFa4ZaDZk7rQMlAKVWXu5XPEChTjxfzXr9iZw8Qdf1rTNBPLxMWO
LS48BLsmr5GXjy67UEUXHgGbVRrUX2AYtWS9hX1O9CEOcvgQiFyWG7+HS9TBB6SQ2461BLLzDSIm
tHQ82QNlJVtLqGTo0WcNrWtZBNk8qWHaU3vXA5QOlhzZmHw9E/y6jLn511lV/OUgJnhM+VkJUv5u
1GWSh+SGQ7IGzBlp1mAMXXSKsY9cSzVqiU7ytCkCfz7j3DJH5ntdAicnI7krHr+QdHoHVl3cPRNN
NTik7Oj2TIhkPWTVsDBGPqiRUwIeX6/EI9jZpwpEEOFrirGLMXLQlE4bDVag+ARha7L0G1Qn/UwS
ejMGqfZQRAgKydtDRMPe5ZVBcXjxlbFRxDPhda1EEu9YwjoxssFUFYaTKNMkzgd/ILMYuoWISXaK
+L64nS9GUjgI6nDexUaG+DxiNSa9V3et6jDkOQxxrgWcmQBpkk37KtycdmM0jrStFP5wmOsnlJFp
SCGPeuT7Jqp7MdnYaR5o3vKVglmGTbwjVEyEhlWMC2Bbyue7NnT/dyA0LgjQbOF69e2BR2bdmIIP
aBoT0VEoRqavKJW4VVJaM54H1gcMOvTiiwzgnJDFqLa7/UA/7wMiCGu4uBnB3/kQzacm2hlKuJQf
T0+vWNMiVBUy2cr3ft0/kuEG36VBq+hWxfKK49u9O1qhxvIIn1z1ZWZZD3MHuAZXojeGQbtv3kru
U3XT+pJVLh5oW7JXXxSWdaz2//oEhs7UgNjE6GxBsIMlGPBbkJ/ycx5yfyxee/gm59BlN6y3qJxe
INbnePJ8joraeLI54HYhmuIWx90XFHYoDJPGQspHtIFbLkbuwDmzVGbD7LA5GRjFnNUrTZfAP1EV
adRX/fDuSPpw1emPPqmQZH5VK30d64GZveWzK9i1yfrdv5e65TEzX6LlxttTYQKkEP+dtczwig//
R1YueNMWN0TwjToe2drBo7oIH3dvjjmCJGzj7L0KVXsa9T9OWhDmY3bFcKwLDrLfrOm4R/IuFEHK
WOdLDSei1hDzy7wy/K8jki8xgNIqCnChyI0UL0h7MGpoJZmBKzpmB21NrbYCdS+XnclyZ4pPkj97
Ylxo6BmW16US+sj65NAvt7uBNJHj+3T8wr3qBqSrSQsvZLNHSB5/u+5ZrPQSNqbhhjQv0NxUm8rW
8mlir3nvxXFJPZ3K+S6GI2Qwnf2OY2Rw6oMPtCsWx/sQiTfPQtb0pb9mnbOcVNeiEbHXgFZ0MLGz
HSxuKW1kexbxYUG3eu6vL1dlUHRKIQ/2irLYTwymVewOAwSODl+75/uB8Wo0kVVvpXGw/mTINAYu
7qVxHRYXpj/ksW4pfMUjP/9kM80OPdcSc/1g9yUPA2RX7QkGwH4JCwwFsIgv1mvu601jFz0O9Bkl
0PpkocFdGAcJZC9DhmjGWZD2cCN9j8QnvkQzeLUERyt2rqFfavwGkaLpxkfrv6OpLM+hpop9o/W7
f/p/JrT5qiANXTGmqz3ylmPoU7Tu4TIZURP/95dqi3BHf6QvnUPTKGAl4uafN0PLzeEkjspNN5/C
vni04/K/QKDpgxa85gtsasDqyIKmwUwKZM9db8gdA4mIUc8FLdgw9dfgKKI4tgB5EpPMO/Tj4lis
tqjm7rIoMX1dCl02nm+cc00Ed2SnpCSRajJwqkmgz9Uw6BQK5BquKLHcV+uKhZLq96f6F7NxXbnC
VSmpjLjMAEWoUhzZfYGWzNZOcaJaQoYR9IXGrPsoNr30J2p3o8wNrqGikw9KYNxK2WvLCY9Mm7xZ
ANoDsp+v7SBkr8eLvaW46it+Y7rYG5klsRcSUw2nGHzcpwmn6qcJp532CjFhZ8hmxQdCEJZIwILp
uVzRdxU2t90fe9mLoXkrhCopSuvSplsAbKZ6yaOhsSOu4PuU5VUVh/u6OF/PfBHMdXgwxU8FGb0y
hUR83gXciXE6dREXeQKuXfCaGYRt3sEnSdXhFFTMqzCvmb7EX97OWDNl2ogFkF1eh8vEFp0cO/9x
ayCzUdCED5U4SZwamqb/MDo9zUz0PLFfyfocYTFS3vlN2VJ3g9+6zxksTm1dsSso6oHVH8ZJP6wd
KIr9m8QKTd0FXZnWiH8hJg6E73Ssrjj1b7gwI40w3m+jM0O4LqBgHZctjoM+4eYsfe85yhVIUyKV
Urgl0O4NuR1uZsW1VMGVtyngNkI31gbHIWv572fxN4ikoANmSxhGNAG8/qCWyXdQfJUNELlRqqQa
kAwhWwDVJZ+k50DJZTz8jARz55BNIjVR8ErTF/GuvisBZVjiueUM3GW1QUQeP/jr86MB0LIYNccP
7DHwyT47vp2fhU7IuvD8FiP6/DegR7eAvpv3T+B+xcT/I0uB2x8fDgPJw1/b7F5HfvZCIbNb5SVH
Tw7kBYyOuTrwFrANCDbsV1429WaRXUdBnqS4UbNEGIFXNSPuHpR13Ge402Mxb5MyuIoWP6pRx+Eg
Pj+pw3+oMLd+I+j8zxN+qdK0FuoI6nIHh8NDD61SHNGXSOeWuJ2wEGqziBE6o/rm7lnw/bQdqxSR
YV5Byzql8lSKdW32uiMMYz5nKDMtqxStIVSJkUCxjUlJ0mnGjcnXo5P7leZKY58LPiS94oXhcC1O
kzKxrKVJznqpGM6Eln8v0BX2ilCKY/b4oLhLU3B0u+qFUU2olYnVfQhZM3E1Tp5gS54P2pdf1v7c
KMuRwNntpy+X5hZYMgazx7Dov2KLO0FXoYNaiIj/o15wKmxexJw2MwilFA9cGzvh4CMHx38XNzKc
wbmBHeWpHQ2ARcOylDwPaiSrZ5E5d47fg7raWfP4ysjybfrEWn85I6dCXk6w0qhPvAXOiW4AZ3bh
xgXiJsP7o766J5nn7rYPh42eWEfuBRnR8dh4lgEAHrSM0gB69R5KiLHVQ5/R4XG1QSCw4SsV5Wuo
ths/6EB8J3AY3AfdjIkHCCeVbt5x8c4K68sXKhTR+ifR5K+G5ToxIAY+OhoJ54flErjCOsmF/Wiu
rfX2Wa8sXm4npR8kPiC5at4zYcE4qRzc0xiEcXBo9v8uBV1Vifu6gh4z5HlYIFA5dGnrDkzIlSIK
dYpVB9FND7PXET8E0tDhT3Flaubox2Hq5oXdATN8WCNhrjM4V/hELCobdz326sZQhR5GUkDcApny
8Tu4F2YAlvhn2A8Ni4Rj3USuxSiyNiEg1PAK3+1XmtcJjKSIl4wJRNu3+Jr2xP+LlOpkl124rb6J
Je/Gg5bnxJndk1c/DuCX3w7v8cZrwLv1uAZ/6bzHmHGswjZVzzR1xNmjDtRzChlCNkuAEz2kRbLx
TGi4H0rYWZ6AR8ZksqJiY4ufxrQg6Ldr8WBUJmMvtPmytfptUDr2j2sHyxEQFfzzya/rhjL11VKL
N7QNG5cVC5N31XO+mpdD6mn8gvddDzOl/qRc6SuOJsMjfPTbzBexpAWrLA9YSaGy/2R7d9hDZvWH
f5qEB1TRWgjyyKuu3LEVeIMTJgnHmeCOujSjgPByFLXLpFVmjFDrB5Aq8cu3WtWI/NfA7Qem5gy2
xsEwm5qpaMi/nT+K4rQPJ1N4gMikPiIoIGI1I9NSxhJrh3PeUJNOh4qrXWU1Wu/XMKwZnPCe9pak
HvHKNuIrD/jHS7WIas9/1iLRBIonDsenldC2bBC28pf5z3WzOe0WPpYYaGQ827RaH73ls9i955f7
qkA82W14/tV1nEVK5kYtL2JaPDbUU6Mfq7liEafhvOXdTnHAKAykh9k7HNAniy5DUH0nnOe3lVjG
yr29Ha3farSkRstToaPVDiM+kHJ8N+TCwK72uI7LbeS2+2LQRlVmYo4X8PY/ASciygc1olGkqFh/
qMNFN6cO7zZhDXiCSeSPwyvjeZXiiGBoH4a2w8IBU2AX7tG5MDMkudV+spTesytgJcAiQs6CpfwF
XsaGajW8R6h291d3smw/AY5JVSjZsYTSvsjofb2Zxm5nd5iL3iWJXoeWWi+3mZQGkXW2BMHF2CVS
71igJE+ptLEY45GJad81yapgU4axkimT3BMSoPqNfhxO5OV3Ta3odZgdYhdqnP+teV2RG/M2Hd/H
E288O8tfTHu90FcsNy/SgvOzLmoPcd0/jHLd56BDI4zowvJ69W1PZyNi2AgFDDHSY64wVDAD0Cnc
6nomSA019TnER/cjplfR/my3/bQV5gcWPTh84/J5wculwphZJOuhElTGmOEhV1jeyaq1Fd1hzTTs
lDb6D1sOMQmeA+lhr8nVt4CThr6LEBDzR0DwrW6HQCfElBCaWqCbnWiKiR4gJSIGEzIn1YHKLcCu
LfEe57KAA1/tUdDDJawHF9BsHlIPOdLTLTORxyTMSOspPtX9NVSGGUWnVvU8FmTNgyVplcWAXUIT
ee9Yg1GI27KLGOkDIezcY4sXmfonRF7zo82INxyaGwCGcRsv8J0VnEuBiejsOBoyo/8OrBH107B+
4mAc3+SyCipuEv1GGPGUbQSbUFhd8bAFZSgTVO223XsnTnv5ewREPpjR9QrBsdWdEKtHRSxfwqbM
mtPlrN3vUor4eQP8Db4NpsWWkzKRD0rVDSpXhpK9d7HGXIHpk4SXGSM9nTh2+e8N/SFKI9vr5mx8
NwwnSy4d0+wgkNtmxRUXUa3IiPFHU/+hE3CDn/4ntwb2GlKBRD6Ae6Y1ehUydDMTz38WN6cs7mwv
juVogt75j5Nk8CmgaQMwbkVFALve36moW/zZokz4L7mitltlw0/FYgtIAe3hqBryx2rQvWDf0C2W
Oh4lru29HTO/+aYwUubowRlHDa0/8At1XdjjdkOuy8rdPtGqpI0CZAJ7/DqNlAPa0gSfKT5Au7kP
YjYpg+Od05YDKTRHtEL8KTagsyy1mcf6P7W+75CEdG4k99e3J2UIXN59F75xz37cnfNt2zwWo8zU
slA09I2lTSE/zMRFXLwpUL2OZTCm8sTOfJaF59d767021lvzPdEnJkGrV2e0U4rQht4rm6Nx7NfE
Ki7tT5Rhe7FyvdRAxRhjmY1/2771QDsWk5mnuOrc4cZz63aJ/cxz1d4UJNa7TDqO2Zinpr3SbAyb
6HYsI3502PxmvK5mWOxRhmbtA5dcuDOFHSCvJkJn1Fim185yR3CbSqJ9mnavtlCY+W+hHZSUVg8P
syLhpJ0i/j2nTpJ39m3cYrFYGqRiBRf3ZDHOn3VFxfWqXpo8WCpeh2cm2yAL6Q6FBMulgN5Z9gAt
oEvw9gP+CTbAiLK4q84JfvUWssnxx49+USxDBjb0IlqWNFGpzv/JQE1jhgELytU0IsPHKFXXug8G
TXYg8h/HyNAKbpnhDyWmCJTS3Z5AfwHCFT2u0sAhLQaeDVFw2DU+IHWOcnkSfnbHElFir4Hfu7rd
EwOcYOgMs5rDiaiTrZwFkK3CKX/1kyMs3S9IgPKgrsXz4uIHvTMzZ3hQYXTC5Y4H9cvlN2Ax/ZRC
0W85mvpe26738kQ52yzmvf7eqJlgl1cNSNii+RWbbZPbk3VhTri/nlMmnwYMbD5gjWBY33A5gqfO
sBDn+F2O6Q6rk4M5WBHKAFleJJdf5IKSkd59TUsiDZvr1UFZCv9Ppxt9L6ZMPy9644PmqeX5TVzT
YeOGylwSDlWtAImiUHOWL3hxFR3XPBou7REWQHnXkRURf+MCBbhOauPVdHfwNkry3/ByP5JBD3RO
0BbSaWAc1Duqhmfy6me5oniY/6iQg/rrtyJ3ZG3U3qLgExk7tn+qxHRVV7sb84TCUojRsjdo+DSN
gk0uEfGVS320FuP78CH98RhDObVqWkjsjb8HxVbFShRf0wHoXjGIYPvSnKrT9VhN+VQkKCmUF7vP
48eq2mtrbmbOlfdkVMSDgUjuMHKhpN7/X3gKEQRaB8ai+luUtEXTKgF6vvt82XMOTswnQmanMgha
0ENrZ28dHSwgE0Snob5mYlafk1QsBazL9KuWopmgb4WsXVR9HxAkysmOa6QShVfpMXgF/lurt2eK
7zG9GMPp+451cr6BwWxmWtN9F30ZuNN26EV6onk+WCuwniVYsXJu5GJl2eATWA7gT6yNcwlnAW3V
N6qJ5Ce802YxQyYHGqr/Dv9TRswto7rNGkIkpVTE1D4mO7zyr4Vby1s/0806/bme07JVbOUotqbC
SVbJ0/W9m8tcKHd8jguDPJ3Wo2Irur819WuhbS9i1LjzNjsckztEWJKcRuCslVYfcrM8VIH/r43M
WxzbhyP+bCshRy7wEImhKIWowgsqM2NUPjzM5GY9NkDtf36bZmYZjvqyA4iXuAy+I5eQKVykV3GV
nd8rbTqJMumcSCIoB8T4EiRkEdX5b9xSrpBVOHyMv+LYnk59mP+7w8WSeDfjkIGuUPpg115vexWa
3mP3L8c/qh/AAL+/IT48uiO8fyheRJ2IXCSQwe1KgTibe6qeCPLnPWg9OutX7ZOENh3f3C9HOPwc
G/Vdf546gc0Ao4Xg9HiXlbk68HCRbcV8SrazEXi3nomQsiTxjv3ZDOQT3yZREypy3t2lJp39xG5e
x9kMEc5NSczN3Sy11zER1sNG4HxEdMYATQaYUaVp7gctY7aRUFeQLWoWulNSVvS7+GZOeHMkHw5/
yRlZwGc+cbBTXZpE+k88139MNA8KTFjmInQ/pSK4gRsUKnOSChFGfMyVoxV3Z3603dBO+eTDGCIg
sqkfNZAlKZy4ewZ3IDFw1R0HQfctegwFKqK5k+b7qfP8TbB9CPlk2XYNoaQ4PV6fKlUOZY6lDZYZ
DaNuEsxmvI792YipnSqZ+NyjfOyyCpH5DXj09Ol1XKNESmxOzpsXSaHKJxV6Dz50wZl78nfMA4WV
uJnsePvE1g/OGZaDFZX7pPEFBcHzHoQ7wa/lPUlxhTuDYaCkytVl19ZJb74X4yCD5SCY7eLuOZ5J
f0zj7uwPjnLMu402QSr7htXY78j0+MhoC7zi5vUVBeqeXvw7vmsp0zxaghJ+DGJEFei2+ROSKqSy
yWvn3lU+b2GvYmpnTWY6XB2MAHuAriIgJ4ruPQM7vf9Xvmc/GolxsRVr/t6UH4tl+67q5X+Qsr5e
eLBG4eWagKTrZYhLeeIhbsYG1ZuiOGJYVIub4e+StYBVEGtCfLzB/fJAsRESKF982kcbeg0M83t8
3UYhH3o3OE2vQX9ez+NRvo5IQF+wivGT0SK55QeQd/fRktmwSBHxIiB1hQiWy+GPj7hwHJs/SROW
8Ul042DLYuUKLkfgKNnWp6A2QkPGvgTaZI5mD4sU6okw8hErv3KCMrtT/DTepa0vSCzaZkfz1D0n
0/6wdQ0UNam4BKxH2AC8FPyVcbOdzlZNiNLUGjDMMIqoqDAJqK0y4gykOMgBn80S97VestIWSCsn
AFFReSu4bCLu3XlH40qljY6wbCw82dEgX8zInQ285Xyr9H9BnpfC0yYVkuNTu5a8qFNVEpc2FW5N
1xHep8yYN3nWEpc2EKdOzDiKYpOzXlsmrqDY4lgGiQHKvHzYSMzlBUgQzrr/eaKeeBcg7lTkXIS0
uE9xM1Dnxrjz4/NooqxChQyRsqNGIxGnTDEZkkNesW5drt32z6ILExYiTPVzNAMKMkWPxLrz5OZO
/RDWzzMteLKyzGbRrbL0UTJqJ7KzUIFO287TnxLWQhnmk50OZ1mk/ZPWebYjtORDeQ/ksyoAcsT9
FOeAx0Wg/WUpMjUC5rlx+9nQYQ2rVVQ3tPe9GnH/AGm/SFUDvpWQ8MYFua67HgTCbEzWJM9796Yg
xff1U8MwYyGKMajYwTqJCx0LvDlAZtH/s4Bjab0Gb/aRN1kF4mE3tO24yRC0DtRyGX9DV7sx9T5b
5EghNagRvM0iftiYTaeJDEKZ95sx4pV1/ITAzm1qeoZad1ybAiiGeqmAzgDuciavuVP7TtuMYiGj
DqxdbI1ay1UVo/e4DfY1Y4+uu/EtFj9DLXKD1jeEtkYPgzgKIW66JJarx/6BLgZX6ES5CkvhU7ja
B3FWagRY5+/iYjRPL/R47vQq/g33VIn6pTp78y6Ez/uUv+LDfGe1J6TuSdZuvhNgyeU15VnRKIym
Lhnm3qtqfv/angAozu26sbPXYzWb38h4dvZGwUZVD/a23013aRTClLJy+QDiRaxeGgF9bnXh8jfg
RnCAYeW0qRvv2DgVRWKFjUGkJQqRfO+wMd+s+iY38Us+wcTD4qWcdW+SgY+7gvA9R60FA9g2Z1MF
c0XSHj2NKu5vr9ztETZjqGJ46nkpduHBoPL95u7CaHDfeASF6yoWxgLbDswJkfLuPAl96TfeSMFL
8VG+f0VSV1EN/CL92AQqm0n6KczWCu/SLY/8PmY5sOTJMVz0dvRyV+gZBbRSPtixs6eklHCOMSzz
pekeY9VydYZEqQ11cmKULGF5/zNgA51lHjU6rRWOoxTRtveEyLiPz9F9zOfSJElhHH6b1R+MNkX4
WnLs82rY/3I/rY1nTNvTZcvmqGURL1GdHLE/c2WwSmWysp6hoitzNoi9stuE+6IXnuDahIvI/Paj
AjxhUbZ5TxlFZ6RTbaAaE8wn7jrp8wlBb9KVfw8SliiEYExYhdbC7X3zIr4+pR7ZDfxA/sbWx2qg
IjSSJkCcjuhnvzdLHBaQJrN1HmNUHYSQUBL6eolvzAzISiAdRNbDdJEtrYD5xUysTi1SMvSylURB
gWywb9XtPlZMnqMPDgNLpS8iL5zbB/mHbQ8HnYPXgHd2d8ecCLMKVuyR3wrU+sheD6NsAM9E1uL+
w86Z2P1C/UZygh3aAzBFK9/UHMAzM5K1LXxk+Gebn4AyFohrdVamFp/cljywjlrpVqFC+e864pGs
fuC1ghoEq7pMFhUOiiLDLI7tmw91bX51OD9hnarCl2zJmpjwLQ4dIKkexZFNTilP7hI7dw3HxvpS
CmVns1GH6E+t
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FF92Y2BScS1tYCbOJ6nl/yrS9tO5nLdkcinIUmduQUlX/rEFHoa3Ivyk0aB+kXloe21LQE4kGkQ6
Q9+cOvbtZsLXojH8eCz5LSxZZmj1OY0HgImQvBdW/AXKvPSh/8qp2AkQS6z06aDmakr4JM27sgw4
e8FcV4tuRcqkGs7bb5nTeggXj+gCM8w1pZjupaF2huj2/7utBwg2caonPL9QnFqNhJnw1y8cEijm
U2tA1t1pCHmc/cfMmTL1KVw5knK/j+GUCQdryhHqwEoaWgcU/WsJ66DlhJyiBG8LqQzPrvznCBbb
LaJ3ZRAbBz91jljSVrMpulWLCnotPmY5QRPBNQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
cqAgpvQThUsKP1YQSQ4a4I/shkrWufEhsDBDReUcDIwQgy0J3zK8Xf8BMFoFrewCsS2KNDRzQ+ER
jCDGccgdbKH/8jqChdozG61idZWa0ns7506SogoQlXjlqxzJaYEQMyNxDX7Ycmqi2PkN9cXJyFzV
5txS0QofbL3mzPtdA044rsuP1fkQj0yHft0ysK4zktjTKWnJPMDoc1p9qdrOCvbt1ZBLB18dsflT
y4tm2j7ie4QPZbNefa8AuI4j7gxnCkSCkqJB+CSn4ks4ndlDn/a3c79q59d4UozEclqodJLD4obY
Qe0wLjtJvGaBIVSj8HG9RNO8kRI3GFa3bHt0Iw==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=39760)
`pragma protect data_block
GMWtVErQpQVB3QwSqSu3WLxWBruia83TiqFim1P5yokKo29mAgXIYlNizSxbf26Nk9QNVAdbugkY
EOSYgUA35K8EugyZncI1gHVntLXQr+gWyC3ZVaJw3i3eAADymRXVB1gTeGEub/8GwoN3Al4EO1+B
yX50gJK/9i7RntmQ2rKZ/e5tPm3MAD7/716l8sX4zqque4O8TJhN6//xHBn7YXthiJpWktmBNUfR
GZkKbPaU8RTsFZmFZp3jVx3oy/gkabMHIYdc+Vxg/ugdN/QLa3zbECsrbUq7eGpBGdsb5zXFExjo
QjNV/lT2gW4JNlq2t80WtEcIHYPZQoaGVGmFuNpcbe3jHhmLtStpfwkhLlnUWwYZtuBbOeh7ZUHy
RGMnDO2f0mWeNsPbnpVqfPdWQW/N6hmaPQ1aH3gJVSi9kve/QHug2Rj1voRqMVL0YiCRzr4r1T2T
+DpIV3VqH8Rtjm5fD4sQjkCj0vUJ7iMMOqHJG0lPd58C50VMg1K01Tse+ympFOWdcT8+3FROksKS
ajyRiP5tUBVcz3BhbqMnIiT8Ieuersbgt+6y5tHNXQw+M+0J1luJotBdJf11Tfcsgxh4pGU/v0RP
VSWsKUHhvhKU4ymrIOWRIb7xItZzMH4U24SK5KsGcCiWvmaOi1hdY4YS76T+vTUAq7k1PFiHbYU0
WY/Xier4NnTtThn/ngNvox4uK506QyHvG9jRfwRnJGOvFieTanxFEok6KfK7yi0N8iElBJZgn6nV
l42Z3dKfdY39zLbs69edgO3uIGuCePlQA4o2iUO9P5g/o5EYUy/wZzRwRIaPlu47LvnLUs7rN3NK
4WBs36WLI89FJ1lQThnm2r/Ghmh/aFFJjRfrLpH4YpA9F4mH3XwnZEe+ZEx9DgHVNnwKOnQ+g8DH
Bfz+oqxMmnUPWrmpRLmciaQog9eYqbDQ9m1S07fiOSRT3sd5TDtyR8grKVCwLgvmVOzVqHoEvJQk
wb7y/lZZlEeJxXzDNdn3asEo7ezJOd+b79lsO43/C6pOJW9dCUxAPCSLUzDlfbUPA2jk2g4TV1v+
hwLGr4Yswti054OqkoneI9Gtk8OsFYsII40LscSKryjgLRMT2b878MaKV6N0+5NeiF6F2vvmO7bH
sGTZKeY2VPsI21gistDXFA+b2UlgcGAwn9wQY4Rvx74n3ANev+1CzND2YqNuo9+4zRGrQWggrhQo
9bGzP+fwbOB9KWOIkghpgk82x5LM1c9q34vUPOFjo9PjavZOH2+98s+xXjHMxalzJ44Sdtl9C4aq
vYL+LFNfuFrVRgo3F5DuDBRdKu/B4IuGctgqBGe9ZdeVYRsM9dGIWfDe8TGVaMX1Oh3zS7ABc4JM
geBa0i1p/c1lTVpA1zcG3tGYlQ6vKLCcFSMXHebDlJW5jx9DmuvjHo2bfUw0evFGCTbDVDGN83l1
OI+KdMh0v5z5K/LXEwvHRP/wlyZnEzeloSiBeybmdwhvv4L2tfkrSJXB74YaJqXBt3HCePCdwM6d
n0bsteAi1wDdiJuiMMKbw5No6ogqmqhmLqKmn+fcl9F0Fa/kxwDxH/KdFzZFsInDCu8RywEs4O6B
hy+HBCExhKOmuPYPEOJoUZo0767bYZ4ebaQbShNJnwHpMGYiFVdRa2g6G2Q0g0f8f92L82GrIKmF
UpIlvvgLgAU8e23cn6TFTvFcyfvS94+tE5b7dLjMXzOcigTYI4RLDfzRVWYwWCiqsWgXxxOKCz2x
xpiOiGrsOTtCnPRv/qldAcIG5frvOp16Pe65fcvUrerDThKoCqwKf84+ud975cyZYwIvrYvByHDk
S27alxtL8O8lAt1OtNOd2KAPg8aKn5LysuWqrF+UYaT8EULvou1+qQQFJ5nRkzEWL5391SdXj0hX
10Ro6VY+rciRoAqPk0UDA4o+K3+VkAjeFa/6FfgspdRzQQWIV4ibcXzMU2J7WZSYv68JHY/6ncgP
VBe+vVaUp7RMHJONr0s3iZ3LSgGHR2/KSSvi4ZfnW11IFF+VgD6K98msWA2NvVE2fsPhdh75rgoh
820S7siPCtFrAUTmZzwyTrC9EFNwueVrj5Mn1FZHbLHCzgzKVk2rHtm/fPhi3cD4Q6xZB7AmIDIA
6wdo2Es8Ll4rC3MaOfsGCTr3N42aUTqi/qhFVEZ0BuOtEY6CbPszGonG4AXUJT4M1LfbbqA9DvfY
dgnnHHxXxBJqAn4YrZlQK/wDpPQRZ9T+s41uWQv7MXMzqeRDq3PcjNSc/wr67wRQZthdxEDX/ru+
KMiBDjSULUUw2WnTauN3CztY7qh5t+KvqKGhQ3bHjs5hQtOFzPG7pz6UPQ6jmLBnPjhn2C9bXwCi
CgLT0Gx4zoIyRE5G1iPc69wMnAikG9h6MQovFa8XHQxv8ejJVJIKJrjph0X5oEvEKPQhNh3wfXi8
xHOjpuJ4NJ8zLu950Rx/k0iLPqKQY1HkhMP4Ekw019D4rvSpGWM2IZopcZr9+hn4GZlz0jAHj2Df
17vF2FhoEwv0S3pr0pznDa692AygjxZq3Zyw9/+Kr2271L1MkaQDtLyibY26twjAMOB8cwRBDiOh
QBgyrbVL4SWKjMJp/tQsJiY2tykXBQXpCS/x760CCud3Rex/RxB4qid0CPKSHtKUxj2UDm+oFHwa
SV14k/m9C6Wc3FpfIGnB1O0fqBnb/b4zbuDmWMwk8NUEn3EuumazNhFp3yt1xiLgwumy2hh0WIP7
SFDjmgC/sG9if7/rwpfClfRjN+jtpyi6D6sSZBgEFHVeX5NWkKwhGd3cC2feZT3du37rEeNxKw/5
CTfCtaLJabe+wXri2pDCcVP6q5JgdrNZvTQHJTIQB2sfLSb2jeCrN17HUCe+5ofR4NR2+GzAjV4k
gxNvYMsgLoQIRnLMtQloGB1QZllUZaBuIUUwRc03WzvX365togiFd+TcS0KN5s+zOgMA9+YQsd/Q
UWW4TIB9EbVI0e1jwZrVIBlZ/s1hMJRNnib78aXs6+Xuqlygishy7oCSD4/K71gvvg8Lw49DAd5j
8HHTMTk4K7d7qiS3srKDq1Ky53zN1b+U4FDJrbin97J/MVM5WmQ2X5xhNSFtSxFE5+fV6jBOW01c
j3YAGs+o7TWwJlmBrKUnqEZOPGpdu6VEC1LE2iBYEj2SJEDz6CKBm58+mZRa0I+xEhpbCK3kl8ku
Y20mDP9MEOaceLg1wdozUI+j2MZOnSF3uRnBGCUDpZx9HGZe/KO2HqWbO8SDp6QvE0EDTepbMyoE
yZWad4t+q6/CaCaO+Yn8YUNfG7m4xHV/o0O1VQU+06zVS4/ubzNh3u0qr+Yzb2FYRStunD5AppHM
RsPai1sxnxMPLzIUxy/FFoxQnY9Idjx9LmV1XJYQEepIbUxWGOoydCFVLTt5MOAwq/OEfGD5lckS
qs+uoXKnpxENvrCNjtiF8hsxKkeBhYql4607eY8cOLB+X9hR5GNdV78N1muDhS5VxVU3089sSgH2
Tbs70ut2/rTI46FPsxJQmWFvPBuszEG1QoWiTiqYTfN2EkQgIRbmXZ2V0nhtKnL14VunxIyudWXZ
rTWI5X7VGSuad/5CrUgR4YunXzHdh01kE+IoBPYqCaoFtCyx73I2tuC88sQIrVtZs71U1DhUxST2
fK4VEaqMtQ7JQGp9kDcZ0jxbpu+5BEfgI4n2p4SnqxVeTLcFNzJzY9+FI2yg8PejyRK4q7RaAa13
e19gB59wdf4k37lSP4dR2zFMjkNnB6HoiVnRAhnzDfV+HKpKBJVEnYYNqAKLTgQMPki5RF6wc9N4
5sCtvm9WGz+fPn4XWqweHffrhGSGl1glSYt7gP2p6y5GfO4Uta19EAf8aqCKKbKtBiPffjshXn22
gqD+rEqjmJXmO4HuBuXgx+3W1e9TJdR9irGM/FMyCg1g20xsZnxzFwvt6YG9OdLoXTG3SfTU4wMX
cb0jdRPNb0M8JOdefhHkGZF/Frr5vnjbBbBI3Pr8WfK+Xex0U3suIaO+FKihleQlk3mr24Q6sqKc
HhN+/raW5ZHT8cnbihocX1KEjzy3yJla3lNJwhjsAyERNdl0BOlgeQPyFod8jIs/DkKhvEDEwJ7M
0hZZXopIkFny1sU4NYZ5UBv4OIrQl0JkeIL4wqiGQRaurdQS+yp12t1WSvjriIulcXLc1KyYZU9i
yUwlUCahewW6yipUNe6NV7e8Hr3/O4W3qJ5jSOzPQ++nsmjBFpSg6+5Eh7FqysOZP0HNJOnSVHUm
AvbiE9NS6PLV4mPlp+RV7Vv5gGeW0kYOOj/65hMqjOqkpRx7SigbMfdzgmCCRhY/Lo59W8ru4Nm6
Rb6V+Uhoplk50+SIqwpr1X+H/KBeOHUn525YFqGQg7qJ551GRfkG613F4sURcReuTsXqhWFoJQjZ
taKpf8UAZoiP53tHpfvwr9NPWBhyfQOpL0WnLsy9m4OWXd6ASxnjprY1YXK6NIwX38QkwJf5v+EK
Hr1Y0yIq2F1UBqlR/vp7k8B7u/Kcs3Otmgr3syMOvNMVYBuXKGewWdRzzxZhgI6yUmHvMmRqGUja
Fcqddb3ugVOnDzk/w2XNcBHawOzF32So1scUUaHXCOdxUuA6AgTyoZLcYX8N30+BBjhPm9GAHept
Qw/cSMydDvGIV7DuZ+E+ZvQJ86Utn+9UfrtX4Iarq9npscm+H9aNEDkCo9gx5BdHVls111pbhmIG
sIainUbtyQtSDQlIDPyGaBX3f/lLvKvIzwtLi6Do6jX7VZ46xTLhxbh7KihKgDYed9Yv6UavNlRM
m9lIMigpp93JNvZu3Wt+NpnfeooQc/VVumewWPNELFKuDPZ9sdmyBzW/vR/oVYAF1qI3l0JK/3mJ
ceDcQWgBj/r1DveHaiEtwpOE9NaYxbTdx0z7oGW6ZJJYreMTGar5citqnsWLl4WHqaAD+vxY9mHc
TjI6B+MkDkki946CGyIeqvPIVzlKEWPGf3Sqle6tB1PZN4ElLMkG/GgFeC4z9lmPPZyTtnrc7NzC
FcSGJm+t28J10vuuGY9YRt5+9su7GuWrLRjgha8BipT2VyqQgA2D/yPV+I17BxZXt73dfVo4Bmz4
CBKrqW6ESid9/rGn9BOk+KpBAo2iZo4RkZrHrY7Oj50BkXH5hEKpPCzHkH7gQqALsBcFs9H1PSb5
eYR02/Szvr0jqr3wPsxp6/RE+jqxBKxKXophbSybEkEePT48BhrdjAOtFKFDfN4d7q+M4CjWtRH1
E6G+qRmI22daRK29GVucFgHOwlgSk0pT1muFecxrugyB38gC2jBZUe1vSoiztkpijf08QW5mWIeI
Pl3lTIyfYAeywTvaqptUMrCICartQuhG1ev/B1gvL03mtcaoYzaKUuK/RJh2nI+GpxQ7JYxPE/fz
WqZu3aDTZt9M7Ddp6GPEu2NOcZ3/QEvioq/hXGceRFRgZWUxfhqQiC3+0b9tffOI+mhZxrLNPQ5g
muR2ovwTTRh8gblnsRI6lLzwOMYl8vgtNtVuh+z5KL9rUsKkLcbyYlY8Hoxin1WinrMePYAnd3PG
gV2QDAKlbnf2lmTfqlZKko+eUZFYeASKGiNqEJdthkEovA0so2Rgccf9hurbcM+xg2R0ZCAShA83
NBhpcG1tsGiDuTVIe5GnFDrxQ2oHbykv24d/jsKZT5kRZwV9+GsET4+vPoEupEhwGPTZTv12gej2
bYVOkdcQ2ySlteK9A/gHW5MoV3DQ19apb4p1OqbroQysn8t+xgh2Z3eS7vW9NoGWRbeIa6LlIqDl
m4Jml2lzd2g38M3MkLzuUOVK4v37gnaUIP1r62GqBePEau+q7YicBBKTG8cdPSc6Sfcnn+s3chh3
DOdRmqpulf3wv2/1vYc86eI9zjVByJNnOlgJ8qmkMudTDpkG54SOzFSqjeoAaIn4lL6uC4SdgdHT
TXOa07Oxt+1jH++gBkNMY5eEQEnZ2owNFhi2yY4pyVAAj2LbssDelXnvuaYrb/05Td+cxa/zQaVK
QHN4UhOUthXF1LyHUuCuwpW/08O0jIJFdOzx6x+H0Jyr7KoL/yScZH8b/LhrMjHYH9rAGCaf5md2
AMf2W2/SIVJE0AoGJWSs+Iz1I/XWSOqfGqKj1DnY8975h5+mMDYQpA0adoFQPrMGo3PH6diYPiY/
DI5kIqXHxBzxDcMdc41p9ukRdpIVkX3osRPJclgRKXRJ/rJIXJeZ3HRMk9VW5OVFhSwLlbWlz2CU
avIWH2yjIyY8HMPEqM65MZirzUus2ErSau6t9EZjMKQagtWVQLE+9hRYZmQXeU7pSfmMYVmdyTK1
pEIQsHROeTcho+O4E8EUpEioUa9hoVH+iJi4oENEIH6iYaYRE5YiZiqwXSfByUTsSw7C+ls70AeT
4i1nYnz7TVlY/w3MNHGCjGMaBWsFgdHGDWnNQpElZKEuTtbtk3/i13rWwDl7XNZno9Efe9vw4OW2
zqHjjEuUH/Kmtt/Lko/IvOs7vC73v+AyRgjBR6wauS52+QqRK93VAi8V3xk+SWowK79SuJZLsM0W
06oBh24Pzpr7c2OLjiiokxR2SiR802QwEAGJW5QuMAJY4otwO1/KaV31NN8NqYXajXD9ttm7z6xv
N5Qgrlz3PM54JTfL/wbXWsFdpGoZWz6rf+EqQ4VLMbPFYR48O2Wkhds/RSdzJlnjJv2eGoXhaiPI
turilB/6B2aUF7bupHHawFlv03bKrkCaccLLqm8D4eUzPPkWbOU/76/h/4q2uwXtbBSnWIaJz+lF
EaYAp5ROEUpEI2XIAE/bquw+pAuCIHBGaVst1RoUIwpVXmF/j6q+8azsFiCM55fSyJmVlGx+bM25
fXFp87BJKFFSh3R2FF5GyD4WuQyYyE+ZHkPAcRnnLSaAbsayZ2bESG70l3ZnEAANXqjwniiD5PbN
RkcffWQPYqfA1myBaXdqbYP9UA5hYT0gm6i3uG4vSAQ17Fxaop6vcLfKSRdQEkKnR9QcDpWhufPf
A0REooAMLYNr3hVw7wTvSEcIVUcwD+GLQxeMtig2PB4m97uuam1DjQy4xw1S0vwRjWT5/3ryYmJi
9A3s9NAz+qhn8M3TvT7lFneZmXJAbWQjj8wiuSAGPzF2MaTw5wzNS9myzJo/ntUFW5TEBz7vNZ3u
PTAj4CNFOf/w75js8EylCQ+AcSMSx5XzF76R4KoCnOrfgtI/N44GZt0WNnafkVazC6mB7hlzvzBS
enS6O7FqXsAh6r62nmL/k2ZppWYWELKnOToSfShzrSZ0m+MJIaIwU0KJuXKgyNpsdSOwR83gZHe2
/8F+k4wVsl4Z6oVVmtoWszY+ioso46ZClKebW00+PlQKXXI+eB4wqNTrPn1oU40u6rWPY59F3HA9
nqMGK3E/R3+jfMcjlvm+z73kQwe4Pz53x+A+OQRfql7fhFjDugc+TWYwCqlMkdqfprnEKjsv649R
lVlPUL/XoIsKD+rCbVXfn0wBeAhfU/dd9IffaMc9xOMWEze8/xkS3QhtttydBmx1JGzwq+JzSRAS
yOHKEUBozvJ2kdQZooKvoCDQolMhUu9FBWnVwxzVezq941Ag+wWsxKz/kSRnPZy3FcVr3pXuqb6f
dUP9Ph9s4EDWNzp8kfryRiJC6LXhzjS3Mfe7p0/MKQ7kYd0BcLJQjzEO/cmPXFx4/YTYAxE+V/54
/Mt9aitAh9hTq/j/2UEbYnmL/xHNt/UNA+8I708oPL9SppVhbTQiBHkd0K4ERrxkQaz+Y9uHb5md
lxJsoNuJQnpM96srzSgiSDXIBMtblyCu+Vfx2odMX4NnDJXJ4DHKa172uhRgYWw7qhQZqjQCnLvG
MJZd3FLEQx3jilxkAaPfZwK/rFwHoDwvZZbxKFil5HculQ296aoEny9n0QxmoNZNn6rfIwUXMho1
dp1Ks0Qtu+U1B/egldnm7m3/OcQs3ot7azt01fgklCtZXpVwAP2Dn289U3hfDU4XswjTA9PjMMPB
9ux8HXt+aJkwXFW8IMVI0AjQDWlL4QlanAlO2J1zNKA+QsIO+X32BcN2mAzIZePwYxHV1zN36gSr
NKIpkHGs2QHJmLJLCtGk7d/QZ8DwnrAAPImkYtZpP3aI+N3Hx+EeqLpGP9PVA6Hu/CIl4zQh8lnD
myaRLqZX9WVAHqkLRc7l+U49nGf5/Yi4bYAVMSqqcJHRTXnNs6gOiuV7DEXf+521HOKt6r19rp2b
SFg9GiPUhLs2406QyiFe2V42Jg05NVD8QiwLV52uASc11vpB4/CieY3B5ucDZOKMQm9zC+SPtHwu
M24MJ2Ul+84MD7dkdob3vnM81N3ZZMnM3zaRxb1ZI3NefdI5GXfq7FZ/ZZnrqavbJenmNOVPN1tk
u3ESmi9ThrDmAo0nB22+iJZUsUIzrpuu1ftHsYv8mzXZxHjBGbQ9glR/PAKMnj/47vhbj2GnS+Zl
7GERhFBw4KAQX56/JIlugaRYVhjWQ1IYNtvYGTJDMQpOoTr19NowOYWG3jjvUp2BSrx402an4qu7
Uj9C6Ji8ryPaKr96K/z08KJgnGMW8K1AKhE3CVzVYeBd8cjtYRmOhzZ+GhJdG89HX8tqZRKWMfWy
zBxnyWOiKuDauEeKHzTNMo2wDb161K4Jqk0/U6kk0JGnWs9y2ZrZ9cIA1jkd5FZoPdmZqtLVrKT8
sLRSs/wtEO5hYdswTc983IMvELQqxgbyci/PICG09+CWUKFBdA9y4+MXvR7abRvbul6zZc9O6NAf
9dJ2A3aXw690Bb+dOOdDrId2AOUgN1wgHsV17VW9Om/ycExbY2T0ofUtvTdK2uLX9tCYdNHdLMhh
+Hj7KXN3w1yh5MHD7zGuOw68bwvI6x89AaLy5CYzmx6M8m7CD8TWCrGi38iO+UP9hUDnpXGNHAoB
cLzHmpX97axCyTyU98Ty8GLNgVwUpRgfor4ZW4vLlvN0EDHNtYUwY/WMJkiAI4pkWfqLqjaVO2Xw
CH0Hsgv8sSeyIsbt/f8p9hu9154zagcDL7tkhcg+Al6I7t3JuZeg6IeAyogQZVrxf2/7PSAmyy48
wby7xmpaFfhXuO+NSL/NUeyos9UkrPS71a+M2hZ0pKAmu/+le864ucOD8si3AFMt+BJ4TJaT/bOg
RnwhOkqTATENkaLWmdsBB6rddBU46TXVyh3yuypvLs24eVJoWMhwfKM7GLVa722JIXTbCqZtgmNg
ctQa9H4QhiR2/iWtjRCpUkRcaouk/ZG9rg6FAd5AmXI2BUfkySUl3xqlNrS9dnPaMe1WozVIbXWv
HPR+d4WV52pTkGUSTLcA24QWCmQgDjgAJxB7HTUh/7l3hiEdjSfbbKqm7qJU6Njbnz1q03l5JuQc
28/tQPZDMvJkd/CsZxUHx9C+3CwgkKHmHxjwCK4BrvlKTcv93ryUTmL3TK/apxcTZ5Znph5xKhy1
VfqqQZ6bHPv1osieG0nZ8WCd3HK30uq3Bto0a3Jfo2C1PN6cpZHzX+Z9sS/jbI0Uru8ZGBnHQNav
00aJLfGyqxlUZm+xI/awZDbtkBL4U6LkmdJ98+44CUfhfG6sF9wTzSn4hkL5u1IulVCvuHPssw0p
dLWjUjvho3BRG3aaUvX09Jc6aXgwXM/tOXkPh2ttBxyjCQPsNPW8iui2mWrZbXui0oNr5mnOcYKs
UTjQpCE7NylM53bKMono6rngYtgH1w4uwpGEy4BPoAFyTW50O7cH61Z36eGPoY2HYlVEtVPI9nRw
/q7CjyeaT92b6ZehvPUF6iesi510ZFF9K22P+Wbd1vjyvvNzCKFOQDUninGxPRUy/yEe2jOIeYkM
9qE34fpjkmjBeJR++fKQ8R58Yr+Oand/YM2k6LYDRUo7ryoZVPOXENsbM4XgE/bCApvMCCSG5CrL
NsWLKdBXfn4iE6yoSXl3hFrZvUPfq0W1VPQAwpnfSLCyrZj1QWa3nSk72iEz9Bwnf7RAO4A5BCh5
J62jd9ohzkyuMFmTDYa1GXIEKLPtaWQ0aBWowiKeRYVYiEijhAqPA1kpnHzfvQvAbFKqyOJ0jlfQ
nDAO1rW1zlpG5vZBiLCWpmGtr45Lsf1ynQdgSGNtFpGLW8Jf3xPSVtGEf1FtGWyEQhoWtdmxkNuC
J3oTXP+NHpgEd9eDae+axm+I1WX9tVX/uaCIH3FxHQZCWOaVNA4DXFvsoIzxWuwALEzeuNsocDeV
lsKFWIjNJV6J0UeMrJfi9W0UV+seQCRI1tjk8M8ben1Pr6FG9Pye5EV6utknf9pEtgYXOpgV2L2D
qMfbsfZbkADzo7JZ7hMK1AWbfAYnLaKxWmhd5Rk44bdo+IauiWrR3uFjaLGCLhnrmwoAhtGDWPMb
y0ar7+o/UJx3Jb4lg0W7ZnWcV/iOQLZGfE87CE8n03WYhS6AaGAGVUPrkptWdWUvYSuRfL/dHG+R
p6kCI6ON9efAIl+A/6GOJumYsrWvCuXXSb2gJghg+H4iZTGeQUOIeX/FZ8tW8x4/AnxJ6jsM8RxU
F6EHv+AZAH3eMR9Xdp8+X4oWADLXnOek7EjP053IZlFSunW79vMD3xwDd5Gb4XeMlmOkfrK6+bD8
b+/LGqJFzlZ2MumiQiIGdiXxxlC8FP3hKqrLKXBEN4PmJW8FAhwRmyrwgidCwGGONUqiLM7NVOhL
1e444vmIUd9ACZyMepMk5ISUE2Rns5m4WxGu+HBYYc6gnQ43XF940ePpaAd+lzcprz0EFcEr8Qk5
j5xCuDnECqiXLoIQ/EARSAombzjQF4v3VNwAZ22heQvN+tmSCO2mJ/FWAIsRe3C50yculi5aO7tC
CQGUIPbiaMsblBZV/5PC2Eog2WxPcTTun7qagIBFElxVVvHgK0T9jmoBL76l/gG6bB/wvi41sMfO
sLIf7T+/1FWtF9c2WKhON/rvk7gw+iBmbFgAEx/il+VEgEa++Fz7zT6fVmPtalI2zS2IS28HMg16
0m9v29wfza8s8Tv9eKZyF0nKggkA1uWbM3qpCudYaqgrRaFawlB9ElMrQrWdTROtIxAqPMFmQLw/
8n4Lu39PIJsk2BM8yQgPEJ6hSat+38O9zOaLKESQDGOywJiwAs2Xd7AMCN0J05aU2+pJVRmkCLmo
dy/sJITZ+8AeTdJHg/UUx34rOxmMuAY9nIPUtvNwFqsnuMQLuHI4jVEZ7E/D9EdCtkn/ndd2zR0M
eKM4BasLZ70reI/VHvRV2JE4a/iF9ZYq/sUTCjRZ3ouf6xM3mDnZvgLLichGaU0Z7evl0iF2aoOz
bQxCVP1dBM+iJJ+OoGtgLKt9yeDR8cDPbOwWCv9/DCsPoAbwFm98BGg8qFYlxyFn65cduuOYr/0W
oKnj+r9PM2x7K7tzOcmo1+HLxb9/NxeA7WgGnPFvUtprp6ED6x/FIyqi12iTCQTq/u2D+4VwdPMY
UI7U4+wnxs34Az78WZUQaBhk6i5gALRAL2oOdrO2E6WYYULV25GC1+8k/V+SZschwAwyJI81q36Z
6A8rrlbsNYRFIlDntxY3piwjQmjry8hV05z90wRG+t+0M9SLgx/oHywg/LfREdLzq8KKqwrlaDaM
LABrZyY0klBYl+6FZF9Efsn8Q3KCbDjibYs8YUNXiGMH37qtl5TBFky5qnzNG0b8BT3Oc8cEWs4m
xFHbbByvRgxB/9iSD20eLhUGeZ1IDMdv6tIbOMq5nJ/Qt2Ar5sTfGWlyIYVJlRfwiGIaRhLj3qpl
tdunyLWOTP4X3TzuddxlxujBypC6qK2wLrjNZBvmOPMPbTLbosC+13VLBg7OTLcUIrduIN0kO4q5
qUzrLxSYsuT0zDzKJz1rfEQpMJ4bb3OGIBVygTMFKRebZYBIAyyog237AZlj4Jig94qLM5RmMsl8
fj5+tKVudOC7V48wjn4zUbuynAL6KWZW2xVpEZ+ixGo4Av1gFt9gV/tDVoIYt0F/G5Z+iuf74biv
83d2KQ6B3Up2EKMW+k6FIfHidhOehsV5SyVK5flgYVupNcPpheokXJqUtFchgGPfaotInh8jS+VI
BWjCf04ysIXQbaOCuAPZag5F2S7NPMaWo5IvrLrAxxv+e69L6MiGkg3ObadZ54DRUxN+6Kd1ihJJ
4uCly8Jx5y3abu2WuWs9s/34U3GgcIv+MqkI30oHlTSI2HjLGYzN7j/PL2+cMaH0AYN18KNm5YyH
SBXt5sKohspy++sABYehJcLJ1PaBU6N1LqjM6+IRE6sOmbtxE2XzfWQ5gT2glKjgrhQNBTDNygSf
b6YIyw1DAiVKBIYTcWOWYn0bNtdTzXq0EF5jaMthtuJptbObZIdzeaxjVcGvkpmT0StnM7TUdl80
QP6RVTiNh7Qv1+rE732r91N+pkVgvHfRqhe3p9Ebem8q34p4YQjEE62liljgf2LgvbsxJjDTF1Ky
G9KYDfumLPfJmtgegLotzwNjCNJXIgyBlCiHAl1qi+9qzQqc8cnd+zpG9PkKPn9+foPE3afealEe
fnw3y+EOMoFZP5NKK0T1VzANA4whqOP5e7mfZT6LI2QB9+tie+QFLp2y/ldhJueAI3vbzV1Xp0+z
x/S95u5KaRzzSuKTCUNmPMP1ZhnihVmgOTvRRt27WMEwVoSUceTy0ySmH9giFyf268NuC6fGSqPv
FtfxcClkLWMETpoNJ9SAPx61h2RUeFS/HFXgS4N2clmnTwDTntzcNyf946mAqtJQ6HEW9OpGh3pW
6fGTKr2YBZWbJXBPDSvo/+6MlOnljFqvhgu+0xXo+G6qXvbNwbmfpRzrELlmp9za1m/Cnm3Vxf2F
+YRo92TGII1ies1fMfpP6YAEWJ3/kXTgVD8D6UXiZYtcHZasgHfyE1RpFJ18JINo09FHwObrV8gx
GgFPE9v54HyqybXRFNe0Mgf1jrIyfLeuTtg0Ff3zJB+iP6h1HZz1NHdJcqxhrxxi5EUbjqjks4df
qVd4c8Q26Unihc4lwppH5OAB9DZC6glg+02ECfHtWUVCkYJNeKYNOsA9N1RXn/XYkwCK/xom3vO/
phvFGwPqhGk/MNE/4mG0e7E8xCvgFkYa5ZbDig2L1EfpRJ3orGXGcjEWCYsoihdmRSVihyXptmAz
w4zQV8foYy97+CazQS5ur5/k45cUIppf0Kvvl9rEA2P2BZCxMXF00QqyIZUuPAJLj0Me9xamkQtX
oV0Px12ulDoA+WBarlTcrqTvtwebsaXyohzlPkvHv9WMAdEsOwPF/YfUZLWH0j6w54FvAwgEcOmp
R5IbBJSagnEIBoP1ErVnZaoUrUjVjYI93IRIlpVOFSIsMeCsGBGNeaw9HE6sVuaxw1g4mZEpKNKO
qdoqAp0lMXOhMMttdfCLSAkgRO9p8oDWr8ihmqfzVQZ3vYU2/mthTCiqYxSjodHFfu8BzFM45PCz
/mCNOLPH4/vXx8Qx00V0p/2RS6bi9YzkOfFY5rIxxbbBeI1QtR19gK+Ax6kqhKfJOXXsz7Tze4hl
bIrQlntiYtrJI68578c7Qk2tqqP3hO5Ol6T2zG/Ia2Wdva9QwglerEGhZ0wbEP7tFsUFd4ocTFxW
T+gvNABqypQsAnoYqpupQR32I+we8Qg5hCpH9waeF3nvKGoHGYKXKD6vFmjyrAzrMysOTN+VkXy7
LLWGp9vfUzofyRC5fPBiuiI9rVT6+tjcscIvvlRvxUevknmAMKWqXjq8E1B9J/DFdHkcZ5lpvG1Q
KfqUy/t/yP7Qi5+AKE8WFOObRaZg765/L5cAmk/0NtjFAF9vv8rCyReF7Cf7NkCEknONJ4NR67uC
T6mLEveqlKY/f1C2ZziOaUtKuCGGuxaU2pNuRL6ayEwKtNIc4z2inWyPqdyscJ/M/sNEuGmT8zlW
ooWbJg8raQFsYE/VjbCjrFm8Sfkxpo7ZA7QVOtx9qIWakzPsiIOjsKEF2G1qXWOUECxr1IU1JXHO
bFhYZO3rTKAH8q5PsjP7eU35UN7S7RYhlnvSD4ukoeXUNkhBqsnvQQnlbq8SX1aIje9o9JYLf7LO
LBTzlVR6FBL2DjntvQi52OEdMFqGHtS6lKS6ju1tMF4lM+6K+eyi00Zt5HY8HeRKDUYk1XWIcEee
vGoCT85M7aGmXy0OqFZ6sRXbF9gwaWDV9IEZ3hw43JE5DpV98HTq2zYu8aQSnFY8MBvNOznrgx7Q
bCik9GGdfyVTpa3kI0Daj2MzHyNw/41zSNhx8FACXJV8CuaeQIhCb84WB6rSWd4GWVVTCfB9UvYA
JUUqOaqUjdNllgN/2R0FFgmT250CLHKKx57ra6lWEgpKOItuFvuqSlsMhVDmEPWL0qrLokziIXW5
l4EYLcY06/emCNh5ozfMIhPmdzlw/eYeKKgq4GfscSDwQUMGe1IKKbxpVtibWazHPO1VHv/+QuRI
ychRu8Wpqx1CtOcLjJa2qv54QMoZrAYiPIpKQJi2b7ghL6CQ+4CoJAr6EessVsXW0F1tMO16Y/Ht
VWAOD+cP8mrbkCt7ITrRPwZ1tI2gZ8zimH+Kge+OfMZLHtF1yJWzdf9BgMtJFCTAEXwl4PPyBfWC
u1L6bnFTyOpuQkrrhE6lghZjl2hOmRqMMjjkUhvX7YlU/3FUK2jtcDupvfazmvJJFOFDWKGsVoUl
ZBB4+adw3yFJn8QkLhXs/fHgNqCJb6AjiCRzAkVpvCGFoFg35gN/dio45t5nYA09ZZPDpmpPB43M
nUuHo87LJJZzRD06pWxW8q3nQhWs7JWAb8HwcCHjvVP50rBh+UzrKYCWNKNetfBN/rCjZk8twCsS
n9ZB/drp/MnTFmsX93EWzb2FtWX2LBajXF1rE17Lk7LDW/OORC6nfyi3U3qkxKW1qFacXe3TkVii
hR5nVJeBwBeIE1Ca2X1SOFikE4HavZH2GFZC4V/+Sn4iTkAa4RLGhN1qszmOgjtl6RxJokoC8VmL
VWbqwjKx6ciiqelCaT3Se+0mzzZT0XJfJDTXkGcCeL7dZFJ6qMTH3A/00LKl/scat1pgaAkncJUJ
qAPM5O3Jxjywc2DDhbJcv6+iXaRm6o+6lYodG9HizjWQTzPXrgJb1tHM7/6MN7o6jUBvi51Od4Xi
1P9J8lBPefXOq8+xeUW4hh0f8U+RG24fMtoR0BUDbATz8wkBZSby1xZjjhDIKFYcxN7+wRZ6gFZw
ThFi89NIAV1vFE4V4zSTEvRRzUXa6kySsIYrgvu3BT/Lu6vCF0wC/2EDkKfXR4kEW0bK9/xAqcT5
Sy2RGzxiFKbtEqBmWXNIQeY+pt41Zhy502ULmliDY3k4t1IM6UyPublJopZSygTR/Y5wpr0DEssS
a3fIeFc+W/CKW+0bk6HNf+dpW0kAfkUa4cWkZ+WR6G/AQq9hQfdauLDc9f/VQrkd7Z5uOqA55w9k
o0KKYiqjkrfswZzYnnpixFwsh9igqEF7pR+nLtc7TBMzFvNrpZBQIOkTx5TKv2NWZkP0zbc459b1
JzNvyaN00nj5ERoLmYp7sAymme9ECfQWPIIT1CQMIbYpWtEahF9wPEbL0b35J9HPLFddap5EwT+g
sFfte1yaOTMYnXJkfgDT5tBtj+H3v2uez/lsc0r2s5uvkDS+zWuPDiS9K2jF3aFsj9vGLdLqxKor
HvwI9EbkxqI4l8Mfp5SNAFawO/8J9Bi6xqPoosNgeQWRCvNH0pBcknwbrx7ZhfNkS98N6w19Hare
LqVKjDsJTgHUyOiripi0nHm0OHI70TUPBmtLEPu7G+K6ykveV7hQsWcVqmgyyoodP9KGtmXH2qnf
P/e/AYCSroyRPUtphawhd5KhdXW3glJWsHHUhqsRY37/dXgEW+lUtF82YRywCMFOx9BxZmb5Q9ga
KTqWsyP9keEN+ztLnWkvn5oHdlq2SRgHTa8pMFBD8JLtNrJOwAm61OLyCINqoivpj0IcdRZztDSM
TOJ5Fn1kQ1PHrAE82Dw3fbdykpc5Y6B5m1XmKxVnto6qB0vbB2GIKOBImKg0DZ/hmMym3OaoWq+3
ARwltGDQC4UKhwUlxyO1XVQuL5hCCqKN7MgZZOf0XRf3FTsER3XfIELK5+90l74tFYxGRFvSiGdi
Q2gJQP0ECCnFkIkkipuZAafQS4yGMVhKW253p6UBxEx/i6m2RoTkC11dg//1XVl4gY6E4Za5HIDk
jSvZ2wsoP/ZjCnWha25/rSHm5MeLnkAU3Yf/XJWMKG4q5Dnl59TKKlXKgKtRC4x5wgw7FwA/rPS8
OtOklFq+9SOBkvyNbrddelkemy+A6W0XqjSfG7SaUfbfbXNELvEQVpSVw3qyjlpckxQ2CQwVSEO6
uhFd4MisNqrebzmXqlGzaFlAoITeSS1bK/2DagaSmSySs1GY2Rjfx1dr/ZiRXXQZ6x3HU3EPNoob
zO0WHiX4xtzUjKRYH21pV5Sp+TFM+LMh9LTWljAHjZwNFR6vkwNP2nuCQPQxqc64K0e/eCDIDY9C
7h7XDaAXxFwHnLxnvSBKyEskvQjc2rwBfAVZT46KFU4BqMIe9ioDRJ1az+Zf3HHnP63pP9czRt1b
g/s/gELzYTKqgb5MHpMTV82x5BVmp7MQJ0TSwJBDCrEA3bla8f61k66je3QX+Ea0xV1BwWpo7qCQ
HYyY4KOd/yfJAtF4nQdV5+pdtmdmznhIQMj7YazWop+dlv5eQgF0rEkCkelj/Djrt81TLqe4TRM0
LQ9XzmZEECvxeE847EbYZQ64EV6QpbcxMDkHCpOqttKc7IqY+lWrPwT6TDI4UufLII92rDQElLa4
PmSQrUs+3KuDhyG19rfD/OZKJ/7meLtDXgtGa2xOa4K3mvaD17wjlBzQg2T2hONneRvPHjL26Dx9
DtD2GnGxrgSkD7Gdgo3WMhXVsvEpWFGCSKjvhU9YnaniKuW+IyfUGJMdkz9WYdqUPvsW0gBvHnaK
dE5453B3Jg7QTJP/6AduJMRYVQjKhilhnThZ5fIgZNLpE3BMI7Yd1DV+VlHpvAc0hR90+tiQhbcg
BAygrryvP5K7B8z4TRtkCe9oZqyYLJVvW6ZNcLA5hKD8gO65//pv7LBhYTm6nXbIeUR7jtQmvbGB
4GmFGfFFQTjYVZCh8n5rLU5qAp11jHWRDEv7o1JbYGVLIlVxEoAOUepThn/0xlFng5i0ONgzy+OH
xC608r/mGCJq6uhpM7W6od+5ZBaWa0q+6oZ4S8jTjQID2JlVM0TtmX/NQuOpPnvPNuGXON3BNht2
Mgxe4PfEuyon2CqZFOXxHjEamum3W3f0fcJh6Dgua1WExEZh/JoPP4WW3buu3eguWsm5bUCYle1c
kE5zd8IdWz1cZOC+WGl/nBcGrAj3d522Bxnky8DaNn1OD4FbyPxXyA1PTc/ZFG+8K5UW+VcpojFA
+CczaIgjkhxOJxXG4gZR3H3XffFXNl7aMufoe4MbaZVW9/e4MZcpuLrqktnEOdb6PKlXd0G0S1PV
+sGrZCQZZ6dfl9Fl4ysJx4/LNyJvymHDmzVyCTgI8fuLbourma5ursvHGjDopDTd/FXzNCullB6J
Q1M1LthNaOW6crp53SmhFGWKJ8zc6PaaEVHYjgNx86EvhIxkRSF/NbNHZP1Sr85oqIIYm7Uk1/cb
ujTTCc+qcSGWmKtjDm2AHvclFqoWKXoL9xR8HAbFeCSC/LQte09jSUBRSMWiCNmmYwEl+uoksHkl
X3PJrKt56Yr4ijPK+08nN+vrFT45TLRFdQkndZ3K8r8+QHvzrBa2IHFLg3TdsI7qgF6+jWWkPx1V
j2kKU8tIT7nhEEofAhJYwjA7ZYF9TWBd8VCNCmTwbZe0foEUzutf2AXuiSzWQRpdOC597bH63Tzn
XPHritnAMKCZ4yzxB12KOlunl7IDvpLm1rFQwjyCwsLX2UVu9RhQdDcTbOsCjDoRcOg+Sgj5QQ25
kpIr/M2defyHGKBJJnB8FM5P21duTQAAbyYHks7gPxAW9jsJLodpUOy7yITYtOKGyel1YBvuom2k
EEA/pQzGumkwtB+ePsAqh/1OWeKfYwqeYyTXfNOC8eezdRexd+4woL/y+Ikuvm23jb44E6VDO+yX
jAecyzjAtKe8M2BvUpfpQI1sSMgw5T4G68FIThaNdgLbdkhfmMdyvaZIxuA0RXNjZce/Hk+HAnsE
WnBMIwpO5gIcs4ty3Pppq5f+JaPXpByLL8wCPq5deXtj+8c+lIiCoQCHm5h5RAk7QRXoTWQAZOu4
DzNHGt6Zv1VGQyfX79YPR1yaJPc7brpx/Zc8Rv0KpvjIN24bVh8qqvduOsLxtQtYXrSycKH/LIRV
RVikG1fr9VoyW9fo0hhTwDmL3NaWGzc0fV997+4HBfYmwNBSosZQfPKZtwUpRFAFW5LPrkP2wJ8m
TSdniJTEYz0kbrejYOs7hXyDKywUNbUIYSapfNiIHd+dSrftwLeOPpHpSRhvhwnH0RRt/aloNrQh
aOnK8trKtuXmtMXOm5/+j3bHdr2L5tIYd2IDr6AJywCBLcqHu1NWJLByHtJahrDrQotMAIkKmJ3n
OTH8PJAT+mnBiScnXb7Gdis3CdM7o4QNfvJXPqyxNK3WNGpOtgQehely3lUslAC5uczlbQh+1Klf
7jzGF+i7OA9oPkdZh2ms9xhDDjw/d5z01r53HM6lG6hEg3hEcvslTSvYCiJZqNE0OVnZ3Mpe561P
g6UpixS09gR1CMo/zYVrhbiQogTKPZDBA9xR5dvUsmWHOxzjFriGIitiH9qDcGWCNp+R1sxSxX5R
A+SR9boTD6FNIyKk3awpytKdtI43m72qRQ0hNXEQXmqwz9XAYw4ilsWmUh9aryK0UEKm9ESeaM/C
Qh83hztHWBn4twFxbE3BLxaUjt74Ecuqb5nftRu42G2yNO4/NuaedYoD9lFFCtsCY4+pgezkk89I
FbfOvmV4eWJDMwDhUbRFQtggLT51GhEaHTMjnNB9zFvXSW9r20cjNX6qJO5RD25M9+nW8ZHK4U22
wnXvAneKcRbMEIh6edoA2mccVvkzWu3fGqxER1CYtkd8dLxIv1HK0bBa7Xmt/HUIkq+dzPPJnXht
G9h5V3BiJ3xdzlrjGiHyAOn5tlcsbInf5eRiS2w2XBfpuwnHYxaYB872OpncLJmnt4A1sFJyLiv1
tXRiX6lkQy7SjxqhJMTCtqtBulSr+BgpqKCSocD8XpxmtNZsqzPL8/YkJReBPsFFLVzflOL93HZI
r+SFvHauQxGSo7lB7w5ocpuSHWdXmIINj1DEYKTTJ+wlvgOLxLZk8L7N2Ti5HezbGhiG9TolXT5o
NGtkXF4i8849g/TWgKVVlXB2foVXHqDQOXqTFCnfyIJUEmmVOP8ULd+jAaYivU3Gxm54jJJidopg
xZai4emte4KGyt+GOZg+VXW2RT0YVtxdMFmpQe6Chr+E5Z7LKt7e5pKnWNdQaHv2I53b2Tm5RHBB
rGnsqBvCbbJO4oK5b028hT3LRxbXvpyVn5iw67CPSCRncV72euIar4OwFXwkHrKJDSlML7/C0qoJ
aAud7u9+VZTTkSy2VCn1BzlxbFeSrA/4grZwQYet+QlAJxkBA4gwdqVfNBqy6NfNygLSjXrc05d/
9Fiz0huS+ZO9VXkJVbs5p89vuKOKYW3t3b3WKZbYVo+9e4y23OiejEbMpJcTVSy5yI/GzNt5MIor
z8Azj5f7x1SfGm8fuwzrQy6awmkaLF0U0qhkB0K71dkMrm4iGjTb6yYufdrhb51pa6TAOKIIVygm
Ss+fRldsBe/6Zhyq0c8UhV7bNcC63Z0brYP77YjiCCJhEe+75nN2BuHGexVO4Yui8ktx0F3Ky0ts
JZBLweVLqUb+Rz/bxpDxjVuL+/OGMeMt6FUpEZ8yk4g1Xgjljhq8/vzTO3VJx5s2zOBcSJaMC5vK
kPUv9IDgkWB2OmnjBoK6rOr/fIUGGwlblO5x75eGyBUk4lOqCKSr5ZyD76cCoMzkg6wBexRWpP76
IDVfIXkx1ZjcMqjaK+382SfkhBr+FMfPU0rHotk0Fl13o4wShoDmyxNi/F6JaaCRKzpitncsMMA1
s6JP/xI3NSehYiwUKF9fA4dgqALnI/S4T6VEUz7Nm0nDDjg0yYs0i/upTs+eBMbXeI7YWpAvSfPJ
ckrXy7IPQidTIXR+DI6SzTOOFx5SiTUqY+4iWOTJnuFkz5D39pzfyccZoNfp9gJTED3SSiN1IuzH
wp+qIZC7r+jVifci41VvRaB8AJ0ilpr4Yqb85mr2UjnnzNrqj/PiuF0kD/kGiKbs7eaXzPTwWDng
CHdNJhQaNJQp2JEHxdWd8Glvtulouo2unqxjkKpC17KjjYezz17KrWF6xKHcCDaKTes9S641ODLp
yssQkUkIcMC4hs5vAbBWmx+qewLK3/NRDr+GZz5YowxutfJyVg6O0NFhOobD+pRO3ffDwn9maGX1
MkvqpBNptYMYGj16ZRmdayPsTz2MJIPqWEca+EC1yFV3/kS2u38j1LzRRHs35EGvNpxeySMBxu0Z
x+UzifHCjGAeAUvqXWQuT78fgDxhLU5Z72QLg/48eks6VmQ6ytR4ni5W+t2hw+uOhKX7V/sC2I9z
4JjgB5dKglhciJHr2lyOqChxRvJbg1vnJZ3jd72KjhzcLw7/X4R3Us7y8ojmO+7RUuAAd4RYhsHk
vFJrX1PrcAh5TP1oYgK32Z4UnFNIkJk3qmnksb+1l0RTyIdTJ1dVD1QfG1QlReFwKy3iCOfI62yO
xTdNhx1PW7RgM87m3v2UTsOOk2ooGMDyv+LSxJqolMX4BCyj1iSoxNvwHD4Q7OkmsWJsYeRY95HW
nrmL/GSHBwH+MtlE4dtL2pdnfaveD46WwhQfSmTJx2+XOYpczH0qLlTi1VB3nkKPlpzmPfRnbj1P
dHXhocRClwtEaLQJrOxWlTZLFqEJTFNCludrxomBvd089OIacPcdbW+thpgBezdqccPOCqh9XwSt
hlm3Koz3IrO6Rcy1I5rVtCaL5As/6S5SlsGjnYy6vKCtmU/SiWsZlmXPILsvypwsgvErZhNa/gvf
NblG1SaAZn2BPTXia7D/QWMXtQ0bnL5wx1xys2XcVZqxiOw1m8Cobu8tBrCo3BSApCrrGJjLSW1c
OMyyPtftAnr3oKYAdt5DJJklMfsqf021oraSeFJni1ahkroZABH/r4QBJ81VTQWixrlOZcBQR/z3
YpZhYh1DH+2eEeKbTp95jeo/Cz/AWqg75lFIzOTSBdbP/xtWxhpR7oAsZKbQzJfl4jXm46G5Ng+K
JbJwUUDDRerLV6yRom5Oks9oQ+ZnEtDwvKqdLXA+floZ1IZ3gkb1tjwtjBK7eCrTyqvOq/QXgzxm
/ewhVooaTqnUV4otAwksxU2gfc3meSCAERVspyJXUqTK2kJ5cBwUKqzyNUqCnEKck0vZPl6KCuUZ
AFovb41n3QB3b2yyEZCARQdy/NYpBH8BiQKbvdgRoYXLgRV2KyEni4FUwGvr5AERq14/DaacNqis
iBwQoQytFYzuIYaeqzcF+Eau0BRsacqXljIS5iRa7JcIf5SNfU70zjgiVqitnXdVDLBB4rsnHtKg
lLKgrKQH7ELJt0llF50clX1cKZ/cY7KCy2pR0daV3W49TejsAv1negf24SvwpEMEX6O6CXsIEiKG
hiz7CbMIu72zR0a3nSL2clkklGlCOjHaFtwoI4go4c0IKnYy9muMB9CFvl8F6LANjcoy1jCL7Bzn
kauUXyq/WtN4+ceTDhnGqsxvIht6QisSHOpwu4NZtFFt6io5OSBqHZy5uDe80Sr6U7yw2gJPxrar
uUvAuXHphGe5zTKssNyNpVwseqjYdxO7Ce+RKB9JPyjtAyJiJ2PxMqoQmHaWN5PI/41uc4tsZvxH
K9EtrIprlQ36QP9Bn/TNQLE1KCi/anL2fPD+WmGlgqjvEVkNKLaOvJE1P7os6//RppNENkkrc3D5
02T/3waxm17Z4DgKD3EKa6+kQ1xIcUFqFDq1Qt8AERwtrziQJ7bpfRq97fVZIlJM290pHDn/iIvn
N2YT9cC6NRVJSdOQQmkE+D2GAGqgRxn5isRc9PM/VjCABUnvEQtvavpIMNVpwiyUpuXwt/CtMMfx
msboYjPuaSe2g+OH+B95T9mzIP9cZ6txzF8gV36g30vNk5WEigRu5i33XCp/1iGJxeehE3EghyIw
ELOjsFSstwzQz9LWa+MJBcE9wK0o7pakZGryVjvR3o8ckG6cJ+vad3qRVTAdujjZ83/bvEuBn8u5
MKCEaUj4q0vUyrQ8JSVDMeoWPxtCiI1JdoM8Ek06zjjYYgGk+6G2U9QC3DlAQ9xWEQNjRV5zYPhR
fzOlRJwvgIqdXVuWaLdPoBlcCWzQPPVAhKf14jChP7HbIdXMzwFMYa5BkrDcFQRqYYWCWEZh0hzR
LJkD+BTu/KAUkHBkkTBSSSPqJkpwKZB7UzgV2XtKHStRcIbGDaB+h10yuBS02kZltqqR8/KFFXYn
QGQ69gsO3ljxTRmJDQX8A/FnsQRCgxsATT53VPbv+nyfGcL0lpsp6cF3IZykqOJ2Mm6r5JGe3hx1
su0aqPkFc5MAGLAErhXt/dUG1c5AUazt3oO6JtgdQ19OKP4YNXcNN20j8QJ55iO5S0Upa1zdMl6c
IBBn9amSF4vQlnVdg56YOArW3J0R/zW8TcBA9krWXgk/rG8jpkwbGnEBfonfC9hyo/5r0h3BeV5n
xB53dtRRhQST78HKNta4LBNrakaXfVu8NvqhBZKFfW96whbW5T8BNqDgz2a+KEjWfCg5ih2BFe+/
lydZM8jkAMimLiOYev/7psw4pHdTjE4CExrsvQtKrJSNSwH1AwgbNVam5bpfhmN5d+pzeO9Cgv9P
SIJfb42QyLgW7nXoNl+3JkXEN3JQ3Rqp4im6Q5iSbw9GYLJ3qNKcpypt4wI1d4anCa04RImXW7pL
Q5ebdbsG5FYpKeQnevNZ5Z54LTsprVdOHi3JJX2jFWfFBbRv2vBLSpXIWmrCj3CKV/vQifw+8HJx
x/rHym7l+ueXRUuFwqj8eek/CkoOsJVLhsb06NbTV2+To8MBQmVlRDSk6/shRzyZ9nxnvwTRpJzH
B3poggQVcycpn+ULZkdxIwbTD5D9KP5r4hrRa/hI9+XsQc7TewpaE9q/QwRJzj/ARnuZMai+bFn+
f1GJKQl35+KA6CaGzm0WEbFtE+abcd7ecixBfX/s3IWYYN4+9tg1pzKXDjjArY9mqOIEGgxm8Wtw
ymosqzFxtQsGsiH5TKJYOPz+z2W8culdU/JwlsLUF6kfw++h3FoIAnlUSyVf4ohaaS7ugh0XLhow
BdD2rdJjNgnBrAkhJZULkcFsTs1LjVOiHGy8xdjocDuEKp09t7HTa9QN3mLzfUxRx/UIRn4IwcLE
oCN2tLn6enbekOStMhF7Veia1AwxmDSz6ch6K82zBWb4IHyTvUPHquVknCWxxr98ZuDoJ8C82kNW
8lbXCKShnZNm5eJ5Yt8jgdDu7vTihf0i/nx/AW2GIg/WK7v14GGAVe9I12E312ZgEKerA+C3ISfs
Y17aM11fqlBqkV4W0THlnluqLX7nY255QIn9skoRfioUQY8OEeerEANi7uSzNTgLiZ20k42BKMXB
8uXnOQRRYKQT1tBtiMZwHEbeEKqiZ3EZFthftxlRLeBqLFUatEM0/fHTCUrC/artkQ6tglPqIIF8
f2VqJWZwrNsdiRARJ3llDVrOE4LUyo4s59zoZydd/cWI4KPzeRnMw8SgG6C3A4bWWWwioFi19UKm
d49hlVsEx27C7W3otg0fAb30KI8hC1WjTz2zeiqVrw61ioAMrFpqfwXCPXQBo0yP4kXMtnLB/Yj2
6zoMr8TSsaHaqfzdzvHlVUTFiTdRVV+H9XQ92jZn/AAN/cBCg+3nX78DL2ShaRB+AZgFUpiaHqPj
jcmfrTblXxNW/lmGdhRaXE0LgEQkdcOWB3E+MmdHzImUf54JAbt76zqJj3TarVobOa/96iumlbGc
QzqYNeTVwYHwMpoJ4Riiwujl3RScH0/jcn1G2/g+VVOT3gx9gGh9l6Y78BG2UU4UTSWgmfoMeSHa
Gmm90GuDIpkYj9gekwTydOntjPIZi6duhs9qCHyA5iVscgp5T+GLHJ0+SMnmxVCYqdb4fmppKH8A
tL9QU5x4u2XD0R7KG+ao/ppIS3fJKLm6AghyHSDNZT84KiJAByGva6WCdWd9h6/71kh8aJbTPncj
np4x4Mz/SJ8g4ujEcS5d4s3nz4MnlWfgk/I09Ny9VqPVDkoJsKectQ1ncncjjG376yZsQEFcizVx
iY7X0rgLWKwyOhL7hxLZ9BVJvJ0qj2fw+sOVIKd6vuwX7xDnrou73gLTpGHd8qoELelB13mGzvnH
MUvgN0R6mAFdAe4N1Nv+mYqP6DSFgBlSiXwhAKtt5N+ZGHpgkbNRnFkeTr8sUHmgT3/412e35/Iq
Wyv7oug+iLGq//k12TFj6a8GLyFF+ACwTjaODxlF88mmD/Fz7GP74MfnrcvJaXSwRwljHI4zbXDS
zMLg2ihNW3420gR9iP0f4VUCP72tOh85rxnGWl88TjrO2Vvq3CZSP79cuLqlph1I/z9ClXxKq7nY
yGe5Qkgb8tJ5NL647eVzR/MO4sEXSF3g/Isa+RKpcCM+7lpCyXWrVlruK9+gKaRQN2UnuXW2CFrY
Uccs+Z2Ggzxdip1mb9a+6311YWPJSgpl3v+lNCOAVJ18jVZYgIZs51/tBudI+PSH5Odyq0xEMqsr
y9paUFYFgW8qUF3QiPzC+ROS3IiXgwI3ztZaqpLwzSeRqxGKvHJN89QhVJlxjc+WV8sZ7wJ91flp
1Kgm7/2hyKnN91PzaXU2j9t2ccoOoso2bn8ygVrkrgpH9CEtJCDfzdvGKghJeXzzHIZPJzxjEpvi
2wICXjjGyqEzuhegfevOuupSdsre/0t4Swbw2Sz1NGKZt/5wgg+VsSfCYpPpuvYBCDJ3Pfqxdr7X
2lK7F6ogpA0E2JacVTQSthvdl5bEnvwbO5GNIfopZvb2dVSYU3lG8TvPbqEjgBBCti+5YmVgRCtG
IgTRw4PG9s9L6Mnn+YeKOFQhR67J2EOvwqWvngmJCsFsLz1wVvC286eQvEzF4MbX8ZZzorlMeY0B
OfY4RWWgtovUjdlkNLsq9G0fxo1wsLE4UH+h4p3YP8CzcN32AmA6UQ+MjXX8xUabnn2bx735tlM8
G2J9MArTuOHA8jMrBvLZKy6NH/Wu76+A1+BVltURbVYU+bPbSs9gvJLk3w9MOZnYM4ezMQlYcD4M
MV70loskbIhZ2EeTVSze5c5uKkBq3poPO/w+biEb6nVQff5vdcqK+byEiKHyRz2+g9AZhdXgZXfx
gfQdKK9Vfyl4N2OjqWX+kxOlDGMhlUIUYEOmQIzZCa0+S/8rOqgek0uTexOpbht0rUeYpj5FZ3zd
zSep+dKQUpYb8aJ3DmXMLtkU7ZiT+xD0uKGvm+oQZlDGgUEy0jIr7bt5oAtNv9YlYKhnnShnsDFI
e9e9PV4Fwozrk+69UVdbnTeKM8uuPfbKANFBzKtNV1sGuNm8RAYXUl6PBknHTNwRKdhtwQzwrmSo
ZDv0tr76Up9WtejIr2mK2NDnDBEx+e+GEjD73RCtn6FC0tRrdcDjkJyEjTUld6Kvj5Aqk7XnWjsy
PLU992BXvMQC3dRIKgsFcHVNxHcxY4zprJv4gEFuHwKuvLrvCimPv06wmbZYbuu5Ct5L95KIIN/F
mmZYRuCvd+madZf+ytCScsaQoo7stjaoE0zJrF9Q+3PeoBesfSE1z4g3d1zudum06vFzCCEaYz6w
UFBUpjaevl7nsVTSss1/86qwR5roWP+GqM7igz6zfvuV3gMbi3RQ9byORr6Dv7s3lNtn0f2A/7zN
oQ4pWuE2lE9ir0pY9PHTC+FcGpznczCw0/SYTUFhapoG0+FpjI23262RGkSn/sctWf1AoPRTsNK5
m6iQPjZXJOqgPpmeGnWxn7QQy7S0xwmA4m4kA+tGbqG/Jc6Zqg/uKoPSBG5XKYv8uiDTf4uFOzER
fdK7Id20y1vPglQmG78qiUMN/q9qHPV4cczTpz0TZJ11R/dcnm2tG8sWjN2P6CDC3FBtPotcWjtj
n0ngot2zSp+Ytq17lSKDXfdtZro6dG51xC8NjVLT0IaolgZKjaVR86cSHm7dnxaam2udhmDI2fP6
DLGw7s4kUtCvjdQnFjK+z1YK9/DhcrXELfemwsWZM4FMYMluMJmG4qjYK8C/Ya0hY2N47ovB1Fra
GNC8h8/Su5JV5ZtnMMVtK1a28mCWcmaxzPuq93JH1sojZZvSlBwh3kjGRO+iCniGfBw1d1KC0yG7
B/aqkH+WXi7Tbv0at1rELlIG5DlxGCUPHtYTo3uyrositvUhqw71UtDWAo9Q8zOXgwJvtKcEJ86o
lrs0Kg6qnFxxw5WdQFgk7jWDLJxq3OAxviFfIZVYjiXNF9Bu8hr3d2Ui9pJY9u0CkgIB4tt37gLV
Dt46nnUpZ363BACkP+2jMHIzDoNGO5w3FeCntpnAAKpUqP559zLU1bIEKvGEZoZqeMhbDSaKDfSM
0J9toC2lifaAsa5wKSKNwGiWTaJfRwtZOsCWVTB3QJKnEytCWgZTa6v0DHEmEPBoYkeH66spebIP
xIpD6Z4CBp2znze2IR3OCTinvJcsTMgd9/bq3sFhJwkKggQH0b6wURuLV1NuGZjzQDCszSh0zZLc
pVEfCxpmCkqpWNiLvF+ksRAraOJZq5/aR4bdibx/CtE0kinIHTr9jjDRwcln5+9mgKuy1GAM94fM
m1GJqihbDsEa8b1J65Y4s8+IyxZ3Iwnu2rY/JHMRpvPCw2sg0tuttL/TFBCBrCn/DxJlPrs7s1i3
In8Lict+Sl+FcDmqCLoHsWB/HHwXgayBmiJbtEvQ4gWWJAVbGRFed2igsinMgNOWyWXOgGe91wvS
HDdbVYg/oVFK/dChKqXiR6MDePgxl6LLFUOseJwuhUS3mAx7HPaah+waiwwt46fy7pPpiL3RJi+b
3K1tEJ57tjw0tH6flnwA/eZ6l8EJTeuKyRq2ry76S17zhollKIt94/IxXLY7wi4mn8LtGLyHJqqL
GtHn48qehOzhyRh2ciKWzjSb46MPFDs2n2TssnDxySTawDzkEJQkhgh0thDvbiZbEmyi4MvPquVv
8IPLjWZBhQ1bBR1zdy34Dik4GNMsWN7Hml/RQj+8ET2bxnyxcN7/fweIon2RMyCMbhuBFmo3sjIa
NQUZ2Q0rWbTMpPLWTiK72TKyJMYIBUsrgcxwsLbnAO28piuHYPdbvKIGQ+EZUYH8fAtTJuI/8KWr
6JZX14UoibkdUv2457tGFBff+oMH304pnUdrEmmV4ZvarmHYm9sF77QtBR5Bs6m1touX6JSVUsAw
X2/P8o9e/PZUThIhdRIYgSvdJMzWvVEFEUYk/ca5YsNLz64T2/ncpT1GNaTvFosBK65Cyk0hCRNO
F9rNdtEryCufuQEyPgA8LFIPnAWOJuC8qcvLGtzxo8wiuVTXeVAE1oMbiUAuZcJW67BUDMoVB3JL
FOXkGJklhUu6JRnYyqppSwnag6nvcjEzSkdKCykIat4AklM6wW7cbqYdUIXkfO6DC0faNlrdg805
vYmpHrNhf2McSdsG66NZiZ26EpnSQ3rDEWo0lSoLDCplqu3upLpL77xUkiVtwAovhFMbq/0qkMS8
2btf/wVthjUmG6bn1qkqvRCi7FKifJ2MNZCr1PnITQLy4mC/IEvlpkW8b17pBrcfd2XdoElq5DBy
hahiJC2MqgTNZSrCIiO0P0pse2/3jsHwz70oyiO60nyYcbPHqoMYXjxFh2GTYz/pzaCvS2l2Vgwv
iRbBBE3xCMcIOBlNISaa4jUe2w6EuNgoPJ2IuxoBy00qkNHsIJirgGVDaSYKlC50PR5shOrq5qIT
RxEvu8EQQrGaxbsOGLMwFUNua1s0bqIIPoYokyzRNrBLN4UxXjWechq9lf0ESTc9i0RCJyzjfZjK
XdsbqWBhfBblUYonV+YEw71XYpz5j6zE7gaW4IAmH700Kgc2EMrxkrxGp6R/M0y67P/KGgj36cGV
q67tWAl4axSsqkmiR27ZRDVyYcR9svbBbq4XACnTsdJNhfyYMG/THST7YCYRKBxbtQKUL0+TRcZI
Atzom5SPZ2+0V8+Lr444IpjKbdzcmMvWINzZTNeQwDHObyWHx716fW4XiOggKBmmnymii1+n4WRV
6j85Du9Zgge8FtZy3PRko2UIdFg/MFk6mt6xWFPHV6+m15Y/NC0Okwam0Syh89Ok8OkfcWXe9PYV
akLR2bqfHPVnUrHlRkZh71k94HQqq9U95v6pCF3m+hiL3dS4RRpDmH5CFZiQOOLbqMkLuJ2slR27
IJwE5GrlchBtsTtZRIE6PBmiTohytht9CGSDMEfYrumL2nwzFdIH3Afm61SJGyhH/bgOq/wZKKLb
6ipIOPstAcHhKbBFM5aoZYofhxWjmodkV+dfmJlL9kRj+ryzC8Pphs+mNoDJu8oWQ4b3tlN7RpkS
6Wudi/9AhYz329wKHEy71iIvIB29ZjqmPZVPMWh9hv1IfOPKJH3ELQl7aKg+USDX/3VMLeFYAZSe
lJRryVYKjQ969xAhbE2I5NxNcS2uR6c8hoZQejBXULf2ye46RUtf+Km47brbcCPi3EIGAa+F7ElF
EJNfnTWG7jDa8wlLG2Qf0sm4HOMTWBIAc6ew3O2J7mtBO5sy391fZdn6K36xdl0VJ6jHNjNRNo1O
8MJDs8wxiVHQyiE+cyChSGd+k7mMIDY4HQryaBo5Y5zfj+l1Wnh/+DFseEf+n+Z/Necv1neFysAg
Z4SWPnUr8B1Z1hm02FxslX0VYqknmIM0MPOHQMA2DDymYPzQb/1hdDHUBdsAgt4zBfZbqgLFayb4
R58DPl5uk0tpXpsHtk7ooQzcTp9EiSOhC2pe0Gnv2JEjQ3JfcPf2DWHwQO6n9/4cUR0JVtLrbMuw
rcaZvOFDVxdZFKqidL9srEBJZBL9O5wH52tfkDU4B7SApQGJVdlafeb71xjiBsFEFVoFvktG5aZC
tlRpBFPOKTX1ZWMBN7luj3u6vJr91/EmpBl+XBbxT6XyYf4OfkvOCZI1gWIKJZEDBUAFJoXpVdAP
//55w9z4ofGVq2xSpiDVEk/oT6gBZNyg+PS2JRgpDeWnmpcJR8NETQDtIgQYhiwuQAqt8tLvKkMy
mMC0G6iqm9mFME46bkJVjY/CdK7wWvi2bmSe920o0Zs8lQLBel9J9AOQnMlUDo/0osiiciD2inEz
VzpmubajAJbZxNGn19UJSM1ZrGASWxdew/3HfllT9JXzLS6NiYveB53yUyeQBzIpsWqM3e7zy4rA
9Z64KWfGVNNT01Ko7xEwmta45X5Rs7Th3HxXH1bfTfCicKr3yrGC905sFBECTbNlekp1J6OQg6A5
0r6D+09qvQYza46oSYDYh/X2CKcmII/waqK32H2qbXlzfFJUJbyP60JqOqvNm+BIoIOiTlMxaKTs
YJe0pez7ETB0jJ7QvTvwDPJBJZKABoSNzH5L8SVM37oYg2YP7FFRRgKEHa56ctJH6k/KE2pALhT/
ntK9i8TpPJGEYl3OEv3fNInZmxh5dlc0UvswO70G/To9WUGILi5Nx81UvxK72mKKEunInwjlr2m8
T+jXCwJKrmdDZxoqgwZT4ZnbpDinzblzkOXrgvvWWZLSIqXrud2r9FM4PxscwKVNTOnE2OKjusmF
n0Bf0+hnkaVmTUs4KsXaEl2/z3LP4xMfhIewrj4hpMJvMnKaLPUyCtnBG5tlxIWyS9UU/31DOTN3
8/WMku0J5O/UnyoCniiioOm4zeLZXOiBQBjPApQA9IcDmmUFcyTPQ89GlX59HGqhlnfyJqSxb54I
TFdYMTomwV8NNEl7QgOPt42i6glTJubsrWtLaOS6tADS1ItGnb60Ui196sZ6uHJH+vXNqWPLjN2n
8YpuZX86lvh8BisJNJSYXxcXwLfa2rfX0hgqI9/76HimoNs7eD923kDVJp/K9IIlmK9ABT91lCWu
c1wqF0ZkBlzarDXTawdpI+QovyqTxmWcrl/MUHWYIus2Cxj9hu6MJeBIsWle6wL8Yj1d761n/YSl
6BxXdfk0DA9rwIHOZKijdGaHTjj+Ra1gZHz4UYYc1Vh3nbhb/84q7phFRMlmxO0oeIWFxlVMO0dK
t35NXJtK9StM+EtdoGQc5FFIz+1RbsJLG/Q7NvW8s8PMq1bhvaJ4O2orI1e3YQm0bPmICIdiI3ag
GMDT8Niu2Ii48ZA8Q7Rk7g+3dTlbtYdxWX60I4uz0zO8dHiJ4KAXz/+wI/4I9ms3WYaTHeYrzxv1
zNWQLO2/fKPPb19l5ocvXf1DgT2ul/3WWvLiIcCfqEH3W2NVHeZsEVA3aHOJCCeMlQ6VJmu+3Do/
CWwpvemKJV+QxOxrnwrA6syCEqxdGNuxWGYeKUiVQ8LNKvOuc2h8iFaX6eZj+6mELA5uRh+RgB5/
8MXwb58eQ4EwKT5/2hgq4mPcaC4pL9SEVe1tN2ksAc+uq5wGOESoH99Qe02bukMsdxGM1K/egLn8
iYzGfQsWHcJtJzYfEqPFOmhyiSoa9jaYMWG2TMRjhOLGFdBUxKFVkw8zqKv+FwaOsCcgmLNrYyo0
egrJSiFEVgYZ3MHLF0dFwWdNaLfPJvM41vGnbzfXiOez98VjFZDO374NiPD5LR4lAeB9GSEdLsbJ
7MRePbhkxp1LiJqmP8YxEScZD/DHLIdizB6pCgn40cgLv2xLQasLO2+2xkl6/7/0sF0EwkAJrHVm
MlNmptjz29UcwhE4oZnLNvF814Lh8rCofX5jKd2McANR7/C56Uc1Q6V96HWpKDxbmZEB3gsKy0D1
aG03NfNIlWEFRNqxi3kk402MbvvED0e5sljyevOe07aJ5SsE2xvCqRjg2euYPd9m8S+rVTE9851e
DJx2WtM4zPpD0wPq/2h4tcDuaYYmfTohSDz1+2CCvmgij0dGNLo1tGaRUbNj8zAaS9HHsmLyG2Ro
HXhWEA96tR2qxHQFoHNl0UMnoXyngQKUCxg9kl4RHzpwEPkGHnXyThO0VPaU+s3e2bo7mSCtARKZ
bLy8eBCwi3rL9kftOadqjAXv+0Sj3OgExjaAageS2kfKJGk1JSdNsVrc9kEJbtm7+oWb/GdDYG3u
41TOPj3neoNIT/fktBXkNXjYX2+QEXg+RmD567FzjIboo9M4d55RfeUtXQhYsfrjHz5qjGDMr4hT
zVdVpXpoTyUksGr8b+93F9dTfk+vPmEUiDOC02gVWAHOXwXIX+Rav0V401rkVpAuz+IAZ2AOMKZZ
cGLepgFEqhxKdY5lBRgr1HBirzkRJd7O0otfn5w/+UEfJAR1ujUIfAoilTxcm+EMHgANbfjkMGRt
HGQbU25THEwHZs1vkXEGjnd4mCi4ZjP1fQoLuUWKvLwn6OkRlfIDE3rfupk3ahg5Dl5/H7V+UKb2
0QGVWP8FYEiShfBYmOq9EDA/yrew5eKeo9SdY8SmuXE8smpZZQDJTeTMCwzFyv7fiEpDYYWuLXkp
uL2rfQW4c5PsjObknWnJrfVfxPUplqoLKZFaZNnMC7Rvz7rzNvklsYcwu0dSsMQsw1Y+rsaT9fXg
SBq4RD2t54wCorg8T78LU+OMMNJ5gT2hhghFK5UAwhvwtZEYsx4VnxacaDxOwF6ddBEJufYzOLL7
8tylpVwOnPVYVbBudh7SqupMzrrVh2TGg28Iivfn1+Z/MgUiCf/b3D1nelUCUoHb6VKllB5+ktYv
M06BftBxzfOE8rESiqxyFCObR3RyaNS+wOF/QBkM/ErdzWBM+jCkv/HDsfj66cnb3+H+sA+CRMqC
1uCTJ7Us/4oGBKZu9zy5ypyfBXjw+/zTXDMd5E+BvQXXl1avJds437aGkugs9/V5ZXWR22g88fob
z5OFaMAgRl3+dbDZ4/rgpb1v6nVdorMawybl3l7WStRyW7EPQ/PnXhwYgVcU7MbD9pcqIrihGVFy
+mwMLnH4kKF7/+DtxJw6V9OHxdOdqGcMiFFpJhpANM3Ux7qNee7R6wyyMAye5rfZrDiFSTewytum
r9CnpRbgIt6UqCdt3uWtMI5UTThoN/vtP4QTaKMAKP3UPW9P2YXmfHNILb4ZUucVN4fVL5LHQirr
MFuEjPqko6YN8HO42+Tjm3Xcq5ImwV12T5uZO/NJk00FRjYm/mqFBNBtIzJJ9tcB8OnrY1Ux6Kmr
R2kCQUrAc9yzAAXa891/p1gOpboCnnTVa7zi3wzQ7o0rqo+LThc3pIc/btn7fLeP5SEp497CTHPg
kV9dUwLsowmbf3CGh5mPx6V6Jol36SU1qCzbuD9ZstNOIebv/sIxcBTs/AY5uRj9uNUYbxQtof/f
pxrfVTESjLJEGGzNZ8pOHA46qOtGqbOR3zaSAbbjHAB1n/zX31GKaLWmeulPa79WeEBpO9sfJVth
mSOqu+QeOys4FmIJHE6NBvIjG7vAwfsdbGSbMYaWmK7s2DVPhRkCLQ43Ud7J3XnZuBh0qXNU/F3J
PV8M5touCWW2yDW0M1nMsJVpQCvdhVepyZ3jBEbC9CmKX4rn051vtII28EPUSOV5G9ioZlDElpTD
LQVy0oOVQQyuYZCaZlNK1BLIVH1uheJduM0RE48YyiySuUyPcdVgeZZpdtR3xJFmLYaaiVTsLPRs
Z83meXWAIOaZH5gRMOWA35jaaVBlAugrKGd10WuqObFprzHxXTvm/49RquPC8OO4kmCBd1Gh2pGk
wYZ3aqc9ifcudaYz6tjtnp6M1WmGCkdFAmnkscVi7GYRUIZSFUQT4jUw8gWNra89vnN1jmeeYKDJ
n2r1Jqx0JmLg992jphIgR0wKo6I+RSGLjadVv28OnL5VXsGxtBqN6QlHL2GJRE/gTeoRUXYeZhb9
2NKyFk96VdR359Qc+i5Qhc2qTYpJoyDffprcgpycmfCZD83qC0CSD7GLcmnamAABXavb92anLEXZ
8ubXnCNuzSQKzxjMrGBwS/Apnx5PRXro/LBbOi41SObZh+VtYxNRlWsuDOc8RCbTGBjnuOy2bua8
IbyBN+wuKYuYkrWeKOiHa7KbCbwcaDnTW/qjWa6mDqeMsfw6pmOjyg9LWIWfwMJQWB4fC6eDKyiy
wJtviBYJIsUOJRqdxSzJ+zn1o4caMMO3n3wi93Niym4e+6qULQm62C/nXGMirJnrJf7fCXuhoUBX
GJaq9vWN88kCBHCn/FdnT4cDeEZKBSawQe2WbU1/wO5ygnI347N4CeKOk32vTWDEiM+NzfYHudNe
zWJ7lB8BSX1hTOxcAPFtJ3tsDlry2Dtfc7G10YYPGRs8ey0+ej9AD13v7InGqoQYXMYnAl8ChI/N
QVCHKO7M2qqI9lIZ0kowVYtyIYHxCteWqgC4043UEZlwH/Gk2ozinjHezcgZc/kRnHM/gMy1Ok0H
ditD3T1qsc13KQFeDoa9Z3Y+Hghqu/gHf3O4xW3WjgEBsqzWUugPdROr8Bg5He8P+2kV0wE5Z5Om
hhn12IyQDHFnE/FWrExKvgzhkxXYYGd7nLz6QHb8/k2Cm88uQknGA15JCzkBAyxe+0/5m/4Hf4tn
5/THBKr5JjvbwR+FGEn/+q4sYkffWcvbxwGcM3TKcJbV7y4VVR2EaR0g95ebxLNLuNftxNJsJUA3
giBAmFD7vdg0a2J2Y2Wr5rc7BZGw95vlpg9aPFtqtI52mml3YWbWTdnpvyVFqvMvl2cgDXZs1LHV
7ijj+g8KPDyY+CnU4CC8GdvRZYYrOsBzUnqcXlneNXqYC4drZnr/f9VsOM7IXmiN170H8UQp1uBO
FzyGAXQ51GMyO3PfX+/l3zbRoHIf677L/ASmNHYrbxL4yh4QiawLX1y3gGZCiPivBx0jKHAnhuy+
Dw06bndIUSq3HC/5iG481siOMZiO/WU7KNaBxpdIAbFnXcQLgh/Ruhw8AqzFJVPwFcSieFRaxGQT
XSXeWrAQQme3yqJFclUKXu0U6qCXG0UoDhoRHa7ik7kNyCs45qGf5qwGA7khjzK6dqm8FFZTd7jv
5YDws7gkz0MVpGpG22wl0wWdvk0afKviGeE09Z0s4ro78APQBQqxDA7kIq6nG9v2gidpB+BdWEm3
J/YsVN7aGrkx+SjhAt3dKXvFFsNIqdBOumIU0i1bWrwM4+8cUboTaUrTpSd3ZLKGEquO5TbSL0kf
DTnEZHKlItamD/fVa0Q9mNrJKg+ePPd56R+zS1zPgj2rkt6HKWHu1RwVxoJ5eMhcoFjSuFxaOTBp
wzMfUhZZYDDR35Iw1orlx8rCPrTIllY1W/qPkKjzcL8UKS8pGg/XQjeTUxkcPqNlD3wzo+ZPrqlN
mkn3sF/Prn6vvxrpeWXjIVtl7uXnppNLNwmxRqVLZQD8pXtL8DLNdHbdLfKSO2PSNblIymXdHyqN
Po07V1yXyeXfhlzEIghT/zFChiJispvIvY4oyTvi++PqptsqiqY5M1xqJnLv+1DCFOmn+0xgxZ99
bJskK/gjPnz52/vbtL18DyZQLFCbSQnIux4Q54VwWgIpDxam4sjPzhM6qx0p4NsPz0AtlAkxyk2+
ZpoZgtMQLhvAGKvMNZp6CqD15896wvGmAdJ2tNQZi273GTH199ZB4WpVarNP5j6TQ+oNKezbynmw
SmNtIFKSTAwGQ6uOOj0ppr9IMVX4QhkG3I5YL+P04XiKTMUDMrYQq81Co8B4hWGNkKaFhZZn0C2e
Oi3m6w7lr9pD21m7GEzhK5seOFUbJ62kT/KAPWTfIyHTnzroCpCt/rPva6UE0qR8HTRlMPYgooJY
yBTDtLc7QPny+tkoF47dvjOe9TH9YmMVgkAJ7I9A/4aFVlz36MGPw4mc9xOCnpzvI09SNcjWLHdx
hnvmL6w+YHnJLWvVT9h7Lnc5yvUstPewCOezSwhyO1YYA+IcNWTpROgDEECiEvKG2R5aruRg7/Gn
GZyd6ZVrt8O3RDecCsKbAcRl/ZwCQbvt1tuYSU35SLma+s2wxiryudide7SrT0bYlfaK0++LD+u/
m/qhdBpEvjR8hJfS8JOfDb/OaU8UDFgPsQ158udCLICJ7wh3rOnh3Gm4+jcHT9JHZ7Tf+WXzYzY9
c9o+828J0AprQS7BKQ2XfR3o1DCNg9Uobmwl4NXLS59nDosYDFWkKKg+CCYpVhBwZxb6EcE7WtCt
DHGFFb770UFk7RrEeohahVIOh+vB9gWauNQgysiYZ66cOipUMsGMc/z+tLtl9xxFiV0Wnaj78HUK
52w/8TENrM5WVyURoKleBWLVpIjCBr26qNxa1gCijn7hzJCNK52KZZousAVVbW/Bo1cOMNpKUcrm
jFqkhk7oNNhUGuLeXd7pK699LJEfBdl8AaiJItIeKGCvmfXr1Zwd3cS/d07w/Hs1CKSDOsEDMCw5
ziZgGUFKUTxlQWCs4hTRkjkhK1SC2hiqI9Km6xFHDAit1ri+ijZVQaFivV3dE9twjnC2To7WlIX/
X4nUiTG3hJ86s09ba0jXx6WD3h0OFkLHizfL/Dy4Ejgl3DnVUgSUI6GY/Cx4ot9NbZOtZw3ccar6
lW+vuXq6PGt8JE33Pi+9e40kDp7jUgtR8A5gzMpa/YekEyP1MNJFbkebj+iI89RYL+lcdX51F+rS
Lpf+J6pR5mK+eLvHBd7pC5IrZ438iUZJo8/YNIVso61yWPqFLlJ7t8xUVgE8Yagj37HXxlYR/zHk
C5wzClM7iwGmVBO5NVLMbOLhnUcEmYDkbvGiGZrS0CtyDRnBkdZi9qEd+dI/xcoa692S4smT7TKb
7eOOHx3+IB7mkgkocT2PQXhjTLR6sBVOBRcVuCmnhxbArSd6lWVBg1xBN5GEo5TaHGiDALYWSSRL
BvcTNyKs8eCovy/SQF+o6ji0WKHv87mdSa7QVvku4k3o16h4TR2lxN7ByC0qb3hvNgSOntPYX+Iq
ZHtAKRJJ7eAUyMawR4irisSUY6aJG1hPGl0CuwpbCyXnLSSezZhRMIvo7NIgJwnePxk35sTKnLo9
+9ZqkbaXEknCaYEcvmYxbO6mTrEjh2FnoPHycpelopUSr/mnqt4YkjNh+Snm8zI6U+B9oH2Enyiv
DlOMhAeHFupbVQQZKnnLcl1x+E69XP5H030zpUPBjng1+hTA0xWCFDkbODkWHlevAZ3f8veS3+ma
Wt82/+mC3DvymY9shznQwObbYseR3cns6uL1anafpSQLsIzZ/pW4z4CtsHBPIqa1OYBbN0zjBK5p
peBeO9rVURc5oCZihuuhWVpvagg0Y85yU7gnVlha0nMGjpHMDLZsIizIOOaYf0+fgP3Opo3K+7nr
TY7tSS/S1UUpufKEUGxDluFBgbz/ScV1/8kzrk3aU+1YpJsLNNx5Tytzg08QtYuqUnhptcje44es
e78g6+kUd5lk2Bl+bZ1srwC+jcm+CwpH3BeR9JabjP2mJeqTPY1atEz3KDLPNsVowFB3CHnKzIXs
JE4SuSCKHMevEkdZbuY1HU54yC2bCFdMeAFBCWNI/HqpVuyCyr/zDvSwbe6mpdOtsmpLQOyzwVzy
d5jGZvt3H5/n20H3Th/HNVfK49h6BU9hy5RiQZHBMLqwG5B/pqpKAIZ2+FFb23z2uXhkTOUmaGDx
4K2Nvl8UiPEWfWljgmsAcUvjss5v7jdR8h5v7nO/qx30pswTIETXDajhGymh+gZrxiU5uujlp1gP
CgrcO5HwzTQLp+nEIixFBgW3rl9nZawXQMnmxAFQwC4c8npPLHeqglegLLAp4ARsCNTykZ+Tnjch
7GHCBMv3k8FRxCALm35ekuVkM5brLwnw/1XjT9Ll6q5UWurTs7LH6XKODnRAdV9a0K/3gOmHvO/+
N37SIybeUtKZ5XXY8WK18ebQLbilzs6WTWeqPbNdPU9fdJka3rlAfhOQQSzU92RE7GGkj+LCSVL3
VrFRwLrzXwlVG4SWTqLMpXxPLMuWIxKqun4lVJSVyX+bEN49eqKcs3QiJbJD14tjhDyQ3592FjLJ
5d7CtxBzJVv6NSLFOlZ/+k3zS+xlaY8RoKH/9x7mKdtX6LSCr/vjYOmR3QyZyTEw+c0MX5Nbjt5J
msKaUxcZGVnzXoJSzPSHL4R57Ix78x8v7ZnjEw2RkwMNih1Q3SPPiYYm7x5kGpHlZpP3+vS0J8SS
EOIKQG+BTmSLaCatxMXn3zqd70cNQHrBlMMjMnBNnjAZCEGF6o+kFAJQ1zahg/+lNNR/O6CXu2WA
HjCNMhKkWiIb4V7IPr0rc7SihWTipxe9crx10M8qKNX5WUyT6BHYClhlD/bohZ35yNSymdEbH1eF
xVW4WPlxHF8HT4uh6jxftrpoP1nZ6PxOrl7tWw4fqVCafAYj24UpCDxCgUTkonqAiPdyt6a23geD
eE3vk3/VJ8kzOpl50cv3hupmfDoB9jjfDq8xghlo5naTL5x1fl1ccLTOebhrSdtLbJwqXNaH5Qdm
Jg0tYvSiYtc+lghp5FRR1bK0/H/e0QdvhdVhB+W0Vl1x0PREUl9AaI73kq9wslTeOvaKX3p+I5kU
TcaqA7WlxODvzf/q8K3Gm0U0EXKtF5fpuV+Jj010SdSctNCzp3MAcO6lPTn1y/uWHYEdIeTIhMgh
+LuENeaaRnvRnGSjLMMzaQPX3dyRmOgoOpsxJ3e1v4+XNbBTEtGYLhBD/4LEAneoJc0WWiQ70eok
AuAUj2rsYnu4gZhZrwKss9936nxMMhYAKhu+KbrypyDaSoYMhoW2h/CmJzkhFZm0+SaM/x9UXAeF
1YS4ZbVsB68mvXtyhzT8vWxXTVQPAaiEcR/hzXd/CvIRG6c06Lvz5sbc2YVzWvHGCPF+jyVbu6Ds
LSdppebhvbHQxlo3MXJ13Mb4fq0CIAuRcDaNA4fNcrQbmYt+B+ITg5x/A6o+M5WerH9D0pP1OvT5
X35Nn2OP2xzCqAynjU1S7N6n2J4rTXnKwXG5jaEw9dnyAXmEkPpxQzNdh2UfBWbhg5GG+yA8mg6W
z23vb0Wsu3I0GVA2PMCxsj3VepvpnLw0Nthn3bjkGU1e4Hdu0azfe/H5fdvU7ViKaztRQFtIFYwX
/yZg4/BPdlfpKaTyfvuS5dwd89omRFhaoQ6Q7BtyvpSG8u9RbUslgtBQ+GMRGsiSKRNGPCQv9ReH
ATU6I8Tm/fhp7WQFf+x8Qg/vMsNDoyooQy+XLusiTV5Q9IY5UMaYT4ZBojdYhLz+cPN4KuXxTMQr
2MTdqwr7mVw9dto2PLZLWuABqtQoUgce0bjPAHDYzL9qN7IOaIGhYSRAG9l00CFUlfBQNsmDzmmW
HEGLIzxF19359HPu9WGcRZbmCT7U5cyMaXfxQlJS3XSFcSEJSg2QbuBQkrJ5Hbo1QN/tHsb238Bq
Bis4FBuxZiBc/B3B8AYt/tZgVg0VDBglG28dq/Eys0ylvOtVpV1ueoReC8ZobCg7Wb2HUDCFK7Bf
pp9Kf81bRuWM4E3XFKUT1SOOua2jHqKt3b5zQY9LLYP0fNTkrKrPN2DwQ9kP6Kd3Vn5lTN3c7hjG
4Zlf6Af1LT80QZYlILnU/iRQAob3QyqzdwGlOgjj4XFfF/n8n1NF3vziLz4JzQnVhhIzMFBMvvX0
myK4c0bh2X7SX4g+iPQlLx+N5DKsc+i0IgeLH18iY95p7RiU67VaqNrColy334RZ7fR8AMtxpOUz
pESRJLT3GhjMSEHiGtm2f3rnSvg2tQItM8nRBlaTv+A4GIVPqNVz8waLQXotzDXF928X3+9pfFkl
F2g/ENMFkap481yrWpu3TUnI5beHX4RNo9MiNfRiitE9VCaKbFVmd+Xn+9+WpwUWi4Z/7G6z9505
xfdeRzI5cs1bfo7rRcVdMLCFsC13ri1XHR2dQPwNIWlSDbWzphA4OoWL8S4//abVkySYZHBD7qGc
ml4Mi8Ay4WO9ES005M9kaYTNk7Xq2iU1pa/IqMxFZ8k7yQDClkEWOA6GAlRNsq5ST1kHdiSMXKJn
W/2csPBfon3unqb6g49bLRgqAj9GtXIxvV0yXJ4BArhrZed2qGo2n/W2zJJStTRohBf8pafFxxHT
e9HnfU4/yS7JeQKLaAT+FJB58XByXa0m4XN0Y0+bjTmmvxg+ooYUKTnFwdaG+Bpzy76uXAfaAI5V
Yk/srCHB6f1kuDI8ERyxNOwyoC1LMf84cAk3qh/zNo7ZmYoPqbvXfAMKOjJoDALIAVLwPLye5uLV
l+3r5y+Gp9AnFJs5oWHXgXBgvao0MNQySgTyCWWjtnJQXaRJgBXLDYItO20xG2Dc/vlRbAX0kugt
q4ZzlwqpqCiUvc2NsfcVU6LoMAAwUdIT0rNZVyZFQJEF2HNRefxZbG21N8UvN2yl0+3HxZzkzuqG
CpqYZa06aBgJBOZsI/YpV/UtZEqL+k/8QMyjn/uSNJUVPMR+9P70e/X0IPPteDHNT/Vftcfwg9mu
KI3B5BsuQQ8yq1zJyf1i7BiaqmzoSFk9UbbNN3OYRaujFVodcWEwlLPp4p1UmMuvcWG85X27FIkZ
ubgcLdGnMP6qZrVeyBiWcFr3L29HIXr7BXdrJ6d0xxIbdqQ3vOi66G9NQXMexbPrBhpQnj3RvomY
WPrkwTSyORzKSsKs62eBHv7XWkEIo8GJiWpRgslgnR/uGPOnYkU05mfpjzDrwhe6u50S8n3fs9Z6
F9QemqTomhRJbUoeANQFAiF7ErM8yu7WaGT9jGi2IbPggDxHXBwE8vgWuIpKKmSdNN0UUwD2JsLP
tBp7i6DcSNpUNJE7DhKuDPO48azmTqdjfbFlC7jLGTtZ4/g0f+BIWVhf1HAywJoU/DELsC22qK2q
mj+umU2Fgg3AWPjc1IkWcjkWMudRkMs4aU8pYM0LWCVv+J9kNZNNjha83Nql1yhUWQQ2QAcKC+mZ
gEQFdacXIyeLlDhb9Yjllam10C9X88Ic2VwhYL2HQ3NFsU6EnJ+Fmxcmpjd9z5FPGB/LaqWj1Y/P
MY24wSn01l6wWfqIH0k76skKgcooRx6Ooh834lYeeVm5zsGyu4jWfuuLeEL1UtH3HOqurrYoSMu+
/wdrcZWKjRmMn4fNf3dpLmSwRG+FilgKyessKU+1RqNA5OeyWuI985/0Vl5KYsmt1sR97kn9UJGy
A38zdZN3Jkb6O93zmJ4Ex7jzGfH8YT//1iH2pWSrRxf49zZJx0h7Wbh3McpmB6j1vNbO78/l26zB
YgVa5jWOHmt8yhYuFkEVq3dJYWrnGNqsppaRYiHiWjp055XZU7Szxo3k87lur88HN5hZhcCwiOve
L/7fI69OC5tie9y67Jpsbq/PvM19Ux16ViIBmSss6u7FAN3Gm6nY0JSKYBHzxmSIwk3HU5fNF3DL
bFYcZ0vYQTxTenGVhBAtTvDR3XYsFrW/GtpyI5j7OkdOAVSUY3wEmgPhhj0p7yhM30LIJ3Fnfznn
3mEEln861UA90X3n8/L9+h2zJAYH9qDwIuHWGcLbOad/uQZ1N2OJOrDwnKH9lk0e0lLghzEpMIiA
GA4wO7+TMxQ/6urnuLwxVB3yU4Q+cpxY+pW9Jk49bkspkhLBog8+RixjCiCJxiWX0dVFGYRZUWhr
xCv6zPac6UnybQZyhB6tPCgUBe5Tge8fAUI6CBbA9ILiM58oz1QdW6V/m5D2R0xPjPAPLe13CJTM
bCkxNasLUMULXM/Me+D7UmUOyIBWKO0nPh9K8LjEHtLnSif5dKgU9fMwKKtmIjt6oPoYt0dLE4mE
h7jH2KCJMowGDH8Zk5kbXsAH9ao9J0wOVi3u718s6LWv+lmPqvZsNXAZhzRcPfO3/GAyq8qOh62T
oKuganprX0QwdKMXgggNj7rm52ISiKAi2CcCKsB/uFPrv1Rzul7KiMyFA2Hcu34WjcgfLG0sh0az
euyZI+9sy9ktkcGORla4Zi+Y0p87UoQJxni69lWZbDInb+QRIlN35OU0DLB4fgkwfVCK/Pvm9dU4
SXKzO6Uvp73gNwD1QUPdO1HW+k1U61WKQZFH5EPHW+AQC0wZUPDvb3aw30uuSONJja1IBCcwxdpz
14VCTpJ0/dVUZ1lY6Q1zNjWkDOxqaFeSePdOa9qmd74XPVs+yX/QDLbcnUgzugegudaezkqc6Wzs
y/8ms8vRk28eF6TfhQv0Hd+yhRNM+z2su9kRE6seAbgfBZRyi6/q8HF09y7BlkigR4ZTGzcKa8Oq
uE6s427WWnJabgs3FEkLFAZkOdL5Fdj+UOR5mu7EMTI5LqsXWFJy3YnYGAOUaZNZ2+lhoEtWht2S
QnA8SpODRbSWwvfC3REmO4CgA2O5R4RoxgDnFPs37/4K4ypFUSn5qRn84ITmSCQzqt60TRY97eAf
yI0unk3fmKe4U66wC74b7jacHeGhuYOhL3DBMwP5XZl7C8KprPumYRj0zPYPxvF5vOGWcSZgk1a8
Uc37ucDoWunmiOKyevXbuIxyUwkethxmZNHiRnR7vYIMq4RPZr1ey10EElzaAEqolrxV7mzw9XHZ
f6cbdRv+H+vFMhqaR1scF0s80yfutPGlttzgNByxvvY8yRy2KHmfq6VfNkSa8LLriXwvfpxFgctH
nvG79Q/nZlX6n7PAgPR0J5LUKGVe5urVclRGWz+nUTHIBoGwgAwUDtTtreWeelnTRzt2TXOru0GE
kHAYX9A3y7fAT+NbqV8TdM1+cC8mG9Gn93KqZbzVeGQbg6YpkRSoaD+DLYpIkOK/Nyx/X6BxHWSP
G6T0kzCHFlDcPLPsjhvp6elmXVoXC8pB/ky0ztB6dv2/WSXBbFRxZTJlXlSQlFiVoG/M+voW+rWK
qjPJBazge1J+l9INPyIjMJuwTeS8ju3e2g+derWlwzxxnJ0ijTtHzONIbIrzq1X1L1uRP7b0fY2n
BasmF54pTdNYsY2G7PkDia/GaBckjUsADBB/IhDsDDP2tqw6YrWvdhN6QHRQ0jewkvqKYDESUwwD
w9SeLlaZA67TEW3ZAQgAw7OF2SZPsJcQ/Waga0Gk6z8sD1mk037gC3CSfSHoVFS+Q3yJ9/oh/LbI
GN9RoXsTveR6PZA9kvGTLEmTdvk441rhK4qXDTu4gYo0EVO8x7MrD8fkUl2ZxVJlX/Pd7nJSQNma
LNFKW7/jTVkpaQpMx+KuZ7tFSeF++9/MbOmFEesACsh85LXbBJPEtWPkOTeJX35P2hQM/2Tv6fHP
gPtat8ZZe2zjA1RbM2gmbSpUx2+qpGLNqNNdvw/H8upnlBj6tLsJSUao1eOh515fKvj4doCIUmHT
eRDowFxSeFYwpC/Q5UvasYuaQ5NkiPhworTmgti5n0SOQ6u+YGXMMGMK6rWpnHYVxxUVOmmgczQx
Iss/YWj9Ml5mK3Ne6p1GIozwz0fSzUzT8LWQkkPTN6LbE3zsnJ71tKav1OXlFq5EUpL2UaLFUZ3/
mcAYbSg/sSLXLnryq9V1xJqPHKFvrJuixFlQ+W+Q2FJSFOAzYgXr9xgCArS5RsSHpngE0e0TM2jR
GVDSGjsIuuJR0tvWoq1cPrQkYgfy1m6Qw47LbT+n2thpDor0l62MxkerDlfBEJKVxZSE2EAeDsFR
7KSyok1OUetHnN+n0KXHY2A4Vmu+igk6Yu7KFbiIMtDUcpvtHiLgDbrVZnxKuoKVcIQBbIPoZBLj
ZjwXlr4Zl45MHaFEQaQ3/P5mtQncnE/0cGStx6Z0yT6+EPRhukz2lHWytbL86rYeBuSa5Mizk3KE
2+3dgyLGkTx1g5h6XBdfKBivH3rRLhYg4YlnJbwtn5PzmuwnEgHMdVJXICA8qTaI3+Q5MUi6uOxu
CKrqOlyACj200ytWSOfT8x7Ayi2tqNpN4TmNupOPA9BSb/ZM7EauUQ+syn307raKGT2oRnmLYn5I
HPLtuko2D1x3B0/bFp3K6kcjQdEJO2RSO/1fHO3IL286UOAXxLTP9RYZ43xIw1h8XC+xUo/5pENt
JZ3QadEwVLs/VMrQP+GJi2fwpIVdY9YsP3RDxcWkFvKVaIa9YLakaZcDjH4oB1p6xdMSBrPpfnek
6TswJNYsoYHma36oNhRp85a9xLbyjs3iI/myxOsPO18fKa0xgp0LZ9+NbyPZLAg+KiFmhtETUcoW
kxuiLxlZZAEQbLS+sZWaaBi23AUkRUq6hhgukKIZoEpOZ+ZbtPXoIwtCZ2SjsW13m3HXCil5H3Yt
97gghoT/1leGFy6CPLV4zs4zrtE0I1DjgQmS6d0dOXc5hSt0LSRxF/giz+l6BEojEVHdvTg/bOwn
3Moef65C7U0RLePyZwYlhYotSB6+hF8+kNVkJfJ4sjKxBcAz8eeusnEplHQgkrPzDodL8KzRgTSN
R/he6UegFPnYEKGfOtx8HDZkxSvClgd1d7IlV2s+Zv9pD3cAWMF74Wqmd9+Db6weFWSqsqQvsE/r
fwjWoUW/6MAaYg7zbvyXjrFljLEo0rnOv5l2RtTtL60PaQ11Wia8USlHsmApmniap5nH/MwxzQYl
KgR0jPAmhfI9mhdUwP7PfKKTafmmjtSggWnIeST7IyVAMdxXRBQtmcZ4t8tOYiS1tQGjdjdHsGbx
xC722nzL/xzPxO+ZoeKof/hCRnunIJ6MFRK+e3H++UHQyIM826DbWcZ5nGL5zEebh8xP/dKH62wD
dJWmb5DJYjGNKTxLG6PwgTZ0K9ehVxRtmGjHEhYNpnGr8jjIq3hfBvkFjEkN3kJT7Lo9Hfds7vQr
eDMDv10HbOvE1T310ixhj9ur3ZfFqCWfpLq55V8GdGLw8ZmT7ENovyVrG0J3yT62v7JJS/LHhWpf
Juqyw2Gh+bK0M2dFBQTEg/B5EfzYca7sZjS8C3HFfFTJWeR0xJAiOpA6iMHVst8fAK6DA7ZZhwyh
jBpgv19cMa7g4PTA8rc9phjyBf7fcPiWACp8E72PhPo1XDyiAoG8rjv5ZTFNb2COm/6MqJ0p94zR
zvrA1CViKbzsPmGtaVdDrsdoKEYx+142TPv4YHQmzJ3f9Ffkh0tVgwEAnPIXHsPRDcfjxtHoGk4/
nEdS+ug2fDwIjwwvP+rnWTEvRod//lD9n5eQX+fz/te2MD8uaMpzeIL6Ml9jc1M0h+Mu6Uti1DYa
9wpjnISeirh68VuS1LYUjrBs5hK/ilFEczjVkUdBaGwes3i9/mvitRkABu3JrpeSsrrPtYoYG6MU
WVbuN2zDGpWvZVQcYEQS3rFL32LfBOSDeDQ3WsfBFQ9/RvzL7chHgBisyndsw3E9erMA0pEQsb9n
XiNHi/brDvle0+8Uu4ME+pHsp6FJu/bQPhLJYa490lCHgoi3fz7UrB1UlJT/2wYBtRhsJvzy6VaM
INqPHT+ZuF+PSuj6XO7zWk6M+T1krANZw9WZz/Xbk6AMLPTrUIif3jv/M+FAcYL3cD+4ZiPyUuTq
WK7ouDugZPKLifaA0fTTNuOoNjDlyv76LBySWdn1tDcXE1jNWnkM+LEhyqicChnGZ+JyA6cjBDpr
TN5CzbWzVACYkozBhTkcOCDOSfq6lQ9/TN8tlqwxpBq/EJ+6lhAl144Fa5Y6BYKSgbXQwd+lCAdI
kxb5EyWVI7I8vJKDeDMnHc8ThLfdM7z1JWWDdwHb/tGPc8Gm5ngKfn1caxNWxDwPhUUm4fRMK0UA
ZWC6YV4h/WfWWD83uzXWclJE+dGVGfu+9BpA6E9mxV/0OLIKXgCNw5F4CJlCkhMllNZuf3AoX+vQ
mAyqG4S5HsLnliOg6BlAsS8+4Oc+pTrd6CWW4mn97qRMzY0swOhbzdLSK3kBwK4V4KMTuwV2++fs
K+38DIpp6bonoGzGrDsmYdv2JVg1edmjBZqBTZtQnUcMOtcFQ8a3k38n0tC4v8t6mTqP6mMAG/8H
Ra9iwM+0/w2b/mnOTqH2x5QHY5MBs8HatJ0Um4Z7NkwI7kSeesgTkPSDN975eyIXtz20bt8bA28J
GOaZFpTkQq3LBzJ+LVlZQK7lvy+3i8IwPo1jt03iEQBjt1QxMG2DpUHvGtSDokSrU4k5Cc/Qh38B
K+yjzs1Tk0bUoon8bWwnPihF94pBa36rx3TKfH2pk9KLcrNMQFeGPA7eTP+ELoBvPm9pOB3il8ew
JsWYiHJRi7PWFmczLxprF/T6hEzzo4z8CZ7RCvTuQU3wD8eyNu6BTvS2saHs9d/68AQxFLxbjCge
7+9XLYxuaNjYntl5MkQG/CQhX734nqlE28sUcsgkYsjrKTfdruSCu4AfisWne1ADE3xbavYtdY0U
GxcXGUXN85NtitIAM3UODp2BvHOm1SywYNyd3WWdNAv2T7nhz6rNcdCP3aC6TM/29pU29QvcFz35
TsFykPZ7nu8aDj3K3HPJYenxLcum+y04f/EdUdkB3FduL+C9DvaZeVDyV8faoqTZkpMvPuSTY3Gr
irECgdNDhY8swbNf8uqH3i/gFtvJmHn719eEkSq9Qt877Updm9cjenzXSJ50kUqEwqk5NxL9h4Xl
FNJsCqf4uffO1+JxRoJjlg1T6J/NBC7KV/cAAnNHEdhLl+W00YmNwToVz5Bm1p/Jf1cBWsJAWxAm
MX5/9ryuclj6luuvAKGotNq1X3nbT056oWw6XMWRUtWFt8/ZGNnWCaL+PAB1uNYbx/QTQ2y2HgnX
ZhQe3s9dX6j5duJRLJQIG9riGriP3RjfoeMtB/X9hRgZ2I3RHANu3taWAGMLBgptUn8lboi0hVEP
9fGnlR84auIQbRLsyp7W7rK1el241Ej/zLWU+ud0oBL6bJ6c4Vbq6PtglzBG1gLeqdLNn+556cv9
gQahjlGH2xKSSghm7Y6hKHiL+RRqPpOBBzarqq3m6iw5ioYa4sqfD7Dn8lyK7ZpnfL8AT5s1sVS1
fsV5funvfrOwlIc30WWIIWc4jo6I+RHBYJDQljK0TDdf2oM2zAIKNPoHZ2HAhNxlkf4M0yMkMQ39
ioFmN1BCrSLQJLQblOiRV2cYiA6gy79MhxzdkuSUK+wOPCcQ+tlLzU31Wn46VXRM80PUXo8rHJ3N
kVQLFFuA30JQ6yacIrMnOpzqqaDOjfVmCwu7GkZonX+dxM03WFofW7nKTl4V7IlGw0Ck1iW1Dvni
VVO4shnTR5JKQeTOqFnfJacjzdybV2vUtXzfd1kiVZ0pTAWLO6HVLrtr+CVhq3dGxFG55dEiQNgI
y8D58xCQRF7T8L2TbJh+6ehUJGMufXiOvZd9FVEMYIXgrhL4IRVi4tDdn86JtZdnQwjqqFWajXFP
BDvMf/AukYDi2BJnpzE6p2Xv8ogh2k+x7FZfL6ZVE3qX9VFtTNRoMjSkGaJwP2LcZehiomxXq74/
JdBbo3n7ghbmSaiHiWc0iDA+KSL9gM/BwXg8nz7VaTjV3I0t1QlLNW3w7Qza+KV4tvQmM62TF7Ms
0Yavc+TYt1iVfdcDW6l2mtT6cghB5/h7zMW6nkYV9ZAvyYQU2ZLfHWpeayqcDXiAATdeNuD/d38q
O+4H6AaNPUJXl12chW+wma0srWIbQfhR3P+F2vmY6UtFqE0ab1Ybp/+OXU2YsLr95ovmme9P+l7n
GD6OoacH2YQVGo4Dk+LtWfiQexbgRXn21T8tgycuNXcbd2v9JbRDJPh32tfTzQOBHyEh8LRA/Q0m
jMojGdSUYPRMTxrrd49vDPDo0Tg4HiFf3Dc8VB6phG9kfuMl/s5x39dZ1USJkqZA0EykpNEAszwR
yo/JqWqq043UHzDQrZbavTENWNNTRXnN5BQrMB5QAaQ8nTuuRucX/26psHBW60+JKT727k9fp6oM
p+O7GfMwOgEcvVc0ersWjTk9T8UOxlf3K20D3ZxKD6WQb5ybKh+cA762D4oZ/T3iw36gyIJrOjYB
yVrO94eT2224H8DUqpRFxB7F5qxjy9GQfcVCtNoY1J91PV9BAbQF5+SCVfm6YArW4m7+Xdd1EegI
c7Cvlwsrbug4yNkoJh7YzpuX2i3WNj+u3kYRqwrDoDKDw5tbKKW8skhxigG82UUClUJy5BrLyXCF
VfuW0ueTALJ6uiH2zy1XQ0R5CD/jAjYbRyTYL7G56McY7ut3umQclaw48JYCy+144lHI7xo+OKn/
YH5+Bk0yReVNOA5Cv8/1LFW+sBr8VStw3B+VQx4DKnYDJJxVqR4sGB2ytWvhhRXiKIIgV0BWwwsw
Kg/IdmfN6tuOtJJ0LiPaGWvdhdFXR8nS/BzFnSCI0EfJ41sdu3gGsX+x5YbzMz98eA8VS5+9GATr
DF7aP6OoHsERMKOjudZ/LNgirTq0vGPsHDw2wwuejY3MVqijheyzC4TceFr3KD/6lZ8WHl5yKmDf
15yqNvuOwKRVzwINpgREKK312Cv9DsisV67BX64Y7Wzzz0aHG3ydFwxLA+On6HlKt4W1EpkEcSC/
rZZsVJqKthxMJbTZpjqgXABuVzOr+CktVqo4P4pea/Ye9JimRGM+YwL0DT3iT0FFzID9D5hO3AW/
HKivWhI5QT4UYI3i5lYvZK13BPW0/6W4QCm28sIRvD2U6Kaml9jpovgVBWH01canEAK7+eS2Am9W
urscLOkhv6yjq2SesA31C+3qoG6PoYQW46nu+7aVBXpDOef1czUSJ5af2sAg79Bu4JUt+L46ASIv
ntdTsU6VctXjL3ClDnASMK0mu4yRMiojvb+KZquh70GA9swAy6bHfC262x7AY6NtVyCI5heEtmIQ
xhnoJOQxybb7NA7TIbtouWg0p9LcDobeerK8oLX4XQfR3uvMtfipIVPgJJk2ZNb7H8ghrXTPPlNa
sKTdsgriTVpqXgWvVwmlBvEjjzOjg5a1otGCa8GTcrROVJiaOiuqPzDldxg5TuOgnnU5ESxCn4mZ
b8nh8ceJika9aiINRTKrH3P+l3flMOg5uwUD49MFeldhZ5J77/HpFLVNzkK/XXXjDnMzQcU2CtU/
/sPRppYkx0/HfV4A2++W0/+CsLL8XmxTSwBL4Lbjq5peiqQTWwsKGWGDrNNGsD+/otjSpwou2lRG
+ayo55uQnhRSHpqt4lLFyawldeaMVNDpUEfF++96e9AMhKkfNLukFZYMebpMJsPS8Zu9q9txK2E9
d31pfjYLNGmKJOW59I5vhkQotomhJylmMeEuX9Gigri7eXem93Jj/J/UsxEDEsUUd7k3GaFAUspF
yZbHpW/oGOt2jCNDe0IVt+KaODSzhFCXNaM42qRDZtsfTtyzPwd49cNX61RU1M06+7rFJ3mZ7LVX
CyIVAQDeCrKnHmqi5Qej23znxLnKY37PxNjI/RQysNvqbjgF3egHSUcNG42kmZJHoD+0Z5UQMVgz
O1neEoZU34QBreqKzTvXuSBhdkw5UHdyAwZmQdvimEQE27f0GVpYnYO80GbhfjXTIn5ao4JFN9wx
rnCq2dIlJqt+nOTH4Bu7W5k2G1oxeoWnRc5KG745C43nm9LkQmxm/Vf3nhkl9VTU7zdAgs6Ev7Ae
/ZuxtE4WtPdpde6JtdXaq+2XNvfVIewHIzsrj+DYY61z5qV6syOKQGw8hlxp/8VJ3THGfrukY/Xx
Zo6FXG9u9c2F5FqCU7vSf4Z/mIZFC7EwTIqsAP0aGdVRIMyo9w6XGH8xGbWq1m5c/bI5xJHzUrlT
ltKctgfHZ9Lk0v3ASN0t1K7EpKUp90kgO3lIUXSThOzCKDHcvwnuXkbLemdF5iZQYHeU2n5sLIf1
TVBKixwWFfKqj53TBOHlLMnbU9DccY8FpZQ8plM8YBKc9+EpEOGnU2XzmfqU7JlofDF+0mLe9Ay3
Ufub3rZPlVqL0npEEEV6q0+xozzrypksLdNQ1GnusqVriV1GT8d7RCOiZIkpzlT3Zmv3A7CxjPwt
Tg7r4wGhafrmfUF4GRyENkpbkbQM73P51yRN6r+GQ5As6qURZZc5Ur6ZhIXM9+U5qT1sdgSIm6PG
XCHuGQaZkPiIfLhQlQ/2+8WQyY6pBJ6PThfwrYDTefwP6jfPb00UgmGnr6AubWkYyWJ+SREbqQLd
1LAzVQVMV4sPAl4br6iw72GNHlTs6ArPrE7Le+yLcJ6Jk5xYpf05L7Mx49mnVC+6U5kECiJpPtPo
eXlAkvF7Yy68q3EErPahLo85B2l6qBrH5+w3GecglzSQw4eK9uFoSys2dCLiSVKi+5PqBe4kahQH
+23XBzgzTjypbeUMiTd2rY5g0FtF0r5GSgoSXnvEnyH53IdkHFMJMSyO3SqxiiXiuXifcokwYUZj
OY7gw8M/BY+23lyt85DwY7teWmYvKVw66fA84ZIkjXxv3icN26bK4M4iZXK5VuoKV7zqL3sBTTNn
SJdk3Ucxls6i5Ud40YshcOhFvEv2fblaBUD27apa/O/W4Y9SFzXczUQFtQusQtqQk1ExOZ1dBUTc
gSHz5XT7U/LzyxrWNzBAwHbEVLYh9+C5z6NSmb9e6kmWjR977/icn7zQWkvzYsLlarx/mu+6eeud
OmpcGgD1YxE+6Jz2B/8UafAJRbkwlHzGe5HnzxKARwoc46a6y1AH92JIGDXY3joJ9mFlmVIujC3z
iWJWs/Zi8muM3xgqOVrECZuIousaDZyPOm3/v5YfMQotkx1Zb4D6RlFx0HMVY/tLmhycRvA6kjUz
9oU9m5nvnOG9wBCQ/F2d9IkMOmJ5udfnypJUL1/fQmzyihcq3xB70gQ5FZ+T4jLdfOalX4UN95qt
tDr8h96FefK+RD+/LRh77sDqDPrFwI++dtEiDF+KFOoozpYxWYo5yQoFgqHMTZWc9Irh/mm66ruw
6mq7A4HxN7pI7xeb/zVzc1+Ve8hLDmD1j6AoD3DTgH/m0r6wIEQqSDVWpfwPSdA/CdZuBpxahF6W
XN8m/UX9aQ3P7nCDdJ9p8VhOLdprwdIE23n/xTB/FbNiTUenvzWNAgMp/mrWPsfU36bPhaKuUe+d
PFZW/jENCkLYdYXMijMdAF6BXr11PeFuDnOVBQHtHGqbpc0ok/+HxZKHlZJwj/phKsNGflNdQS1K
xz7GSmkcCdumV8VRr0Lc86DkaZ7AA9O7vMVZ5/Q5jSSFCZkTXqVVTD4b7utFUpWNilqi3WM86XgS
lLutklzj45sfyYuaC0pbjAiQCz/B72+gk6OR1yG2RNfW2/AYGhybtu1ppmOVrLDwwU7bmBXtI2om
c+rxyh4MkA2h0Vef0W6Tiq/dsluOt5ANPL7Ro7pTDkAUZfJjMeVpht4Xyx/lAhjUfdGrjG+5DTbK
/8YFDnGNSY+wWQL8x5wRUA4ZFFJjuUnZK5xxXn1KkG3C34d0+ARCTgJESXvF+Zb/03vsvlg1Z/zl
1hCgJMtYhdEdtqPNmIi1UDaNBZAHaWKI7vhCP1jlZG84VugI+i5Fdj5ITzKmPG51L+HgVjkV64Sh
48J1sLsqMef3z2zLj+UGePn+fhT5Z2S58Dgk8/VSwaJBamK7g9t70TfAor4K2Oe5Fe9F86QPlUsZ
/Ls15ZSEZUZedSR9lOCvu6z9FTm7bQnn0ugtaKTzvkooarM9L5rd5jF3HdbUMMR+UKUPB2jXc0NI
GZxXfGoVgYHU0CtT5attpBH2dJw80S+dpLyvqJNeMWxivCA9SXpcHsOwzRSGvQAoYdspYIfhPt/b
lz9rbWo0TYvy1MutJIULDVr3xmAETn4tLFKRKSGy5hZzqCTQq3Ke+cgE60xLfhQbzMMlbsg0065U
5K0gTvx9zwAdOK111kKgMU3jO94ZBpZYD2StJdXkoWUWxprl6qOJn8dBMpdW91K+avAeXO1hiEan
a84+1YyhNJIIlLjYDWgu833svV7KkOlNVUHYV5DKxXPoNbYVoTLUdaa+LGVV1rZZlXEBm3C7D3Q+
NZVjQtU8WKYRI9TYDcJW3YfO6eQnl07LbQ8g+8pOtFxdqFTZmwolenOXoxX/j+TuvyW9Dxo1JIVf
FOayw/peEFykHTzVJQiVUtC5ZBkH0jOy+FyCmjYN69YKyjRqSA2jDiXhamzT3ItsujEjhTDKDm7m
Q4mDQ0IKQv33FKlJBBuCRmg/tMPCeac8MNc4DZii49onkqWm+g4J2+CSilLZLQtlZg/odUajXaxh
SvlzqG6z/4mrxKCAmLjTBfygjm404DWkn5bHzkwjKqbrn/35R9nFgp/J03IHSIkDZE2d+W0RlOw2
A5/CPUC2e7WaqRHsYpO2oItQmAYHqiVzbMxJPA+5TGkOkhz94tFECfTgHOwagGq/PCuy8NhadOX5
pLHRrwst+qMy3abJ3w3hjmmUUowQLqL1zMZDwBSdZoXMo+PGZBjqfvOabG6k+CdKCNm5rx41AZmN
/qaF9kJl0tipvf75JQxC9gCNRhWN1sMPieTNmBXPYCKCWZkjk2geOXqNNevkLoArstiLmhfE72Yn
W+/edOH6IYRu8+L6caM5PSeIR2VeE+3pR/VZ2KAEsfaWr+70Kpi5sIGyXCAtnUfrtkp4kT4rfR6/
0RhYwMUbUwhbqSbCsrHQE2ZC1upt2EvFyyEX+whJ/Aj4OmUt7y4EBg0/y4QUOeXJI+xXEN9nYAnw
bc0niEy6ngEPQ253kwY6dKW37Mkcze/QgF3UbbzyWeG5+pTzwcnRC1+6PvGvcG60g9eO3BL20c+F
HJr2HwnWZBJS6xAg8Cm5+HntYK3SbmhEeRwIA2crhj97G07JHZYqczZDc9sTOKrRN0xmt/SNGzYv
ZrO1xrtTFuiPTGQ6NJtAQ1Hdb4CyfTx/FWxC8DerzmCMmSPvDBkT7o21z6CVe/ZsND+cejbGh4PV
dQC4byj5ArzgDw/Bxi23JJhkbbkfOZ6zPH0REHLG2AaHhi8IMs7EejoQxzsWOdbezK4KG+T3We5H
BkpsIduwqlhP59V6NS/mhqC8M+ucpbJkW7PSOuUfMiBS5bBGSXgS4+73T3LPm3CU40IaeVF/E/WC
vdi0hZp7FuqKsG7zDlU0k/8w/t8xJ8emmg/LkDe6asOek6KKr7XrPuI8giYBlWRNpdNC/6Ezkbkj
jefMmd/od5jtmEVmWgq5RUgcj/wRssgZoxvZqTOGgIGXiztk+AEj7OzZAvsxxIf9K3RSgDM6a763
cvg1YOXwppXAr08PPHbESvhKR1byw5KceRZQO+iqBBrSNLqR1mUrqrhNqw+gd30IWvPo8A4gE2tY
umaKjGy9+cpGM1z3+Tosmg933WAaYN0/itkq6qu/PwoTWCf9qOxJ8mBalKDP9xLogdhBxGGNbEbh
vYVyel0xyeLC9n7Yz/6p80lGPeYxlXe1H6qy64Spo1nHBVXhGX/HuNjDwyng+oGlL4tZJ7AFdKoa
OmfLMgSfLQ+uip42G3rdf0kAU0FAfqiFup5/TiPfRcGzoEvfZZynLBV4+uxd3AAE+5guVDVo1LEi
Im0pUoWxr1bsPV/BF2Zy+MQ/zKiZio9h0K72sdO/R1nw3YbMUlrrGlMqFLzUnSkYR2VB/Kh5MvK6
7IFd+22K0qnaF7dVoIdHG0yy7iBVJC5xX/Ob8Hd5QAOiCRtplIHmMAuD5r9NQGvFLq9OT1Vk9ux+
C7gtR3KC6YiAu2V5pUetYcVEyYYdSTl+oemDK1zaB6hmr6AdISeqwW8LfB3CH9x/B6jIctv/ZoEC
R+BjWXb/m5fVK9CFHvpWlww537ZDz1wpC3IVl52lIBDxYRKGEdPMEs/Ll77t/PL4im4fINT2fnIw
A2YaliiRHZeSj45XYExQYfM19ea71YbDfAdPkS/lHI9oBq3o4TkzkinovDaMRA2VxJnseIR/tcwC
ambTdCmxOEmiXfhuaO/QDEztTSYOd/Et2C6IMw+OOZtdRNmgIGOURmKwK1v8StI2lYO7uHhMg7Kb
piOpGQmEvQorZytrqkDOAEWT8cht3tJzGQPBnaSWdyyg9RhBQCwjUXmifq0t5uiZ457LKtbkAx21
4NPl04DOQAMzI6mLi3aapCN+jRsxmmd9bEGPGwK1gdF4DEMX29br3AQEr9TAR7oL7QSX/Ta9H1cO
IEDFHXXaFnwJCVCfLLnKCGW7py9mikN97zxB8bYWObuIh7M0MJtAqa3STa4AHrts7LFIHs3auyT3
r71Phd5A7Uio7pIf3t2Pb0sET315eXGWYcuoG69ttQ==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xI5rRsZ8D/mWscsXgMgqvONi1IR+WUmvlhOeHpoqbkmGbmmCKddy2Qan/TbchxUow2f4O04cfAEu
JYQ5L/DafoWEAHShGyHztGxj4EyJX7x8yqtcAWwgcJlMfy/2Z+sYHVx4ASnUNZeQ8HXpWibYIZuP
FjkTNuAr1SrdQnqwhH5cviaA/5OheQSigRQCP8RRQlRyBxc+biSsCZMpGISZFX2CZjSyU+7V2yWW
ay7r6zDWmMmDZjudTCI4MmCNXIWpp/bhBBuYrBSF+L/5EsYX/jb3bbE7tKSBxKDVS/NsrCqqNgPq
LE6lSb2eW+8BDcfgsBxnkhOXEUv0U/y1UADlGQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
kt+7rNkOSYrcXqbgq36Tjy1mVNbqyEaJJcQomY0hj5jTsV2loT+ykCqTokaSF04RFimKeTBrbOMs
fGmY0J0Y3FLdb9mRm02LfOxlSlD1IAUzPqmK1XSR8d/4MtempkKY0sPLjad2NV3YwFQOuIgbOEwQ
WJexgoWi794m/yDoUFziRVt8L8gAHObe8TsXdCCkIFw1w5BV4qiVphOfsBcAFfGjk1h0eqKL4hHd
+knMywKT44w7gE4DaneMKpcCfQ4X0hNR6jP67PdO/EqqXFjgnAn0wypmmiFT+lBYDb/eP0n/hSzE
W8aox1YjaQtyA9zwXG2XZMpfhHFKcSJlD/u2/Q==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=166304)
`pragma protect data_block
RvX6YNnGq/QfZrX3+SpkwDzMRMPNyB83XtyOs+h+gSiynn1XhUeSuYChhjzO2tVQ1rH3F/vCPrla
hD6VUALEq148nibJmMdYwv3hTk+sBmRcjCK49iKFYZ/tdhMSsIm1BIZrY8EQWICi7teBeErv3NJb
dWXAjbrToZfLhLs8dbOHQ5IeERmI2jxMHlIDLlxjLEHqV9ybINIEoYCUNFIKX8yrNAOSiB62AVk9
F65vgb+GThPHJp1sNpOWimfOv+/6Oo/W6BOOxzOHMKJY1us6t162gsKUU0fWBNrCj+vssOQq7SrB
crH9zn+iMCxEK0YZzuJkmCMWqZ7AZwtfRM+qEZNUA00xy4hADuAOa/xj7enRywhQzcafss6zoYIt
1lhyGaSALH9yhQlAkHYu1D0CdjsF2iZjIP5bXsPkxW9PLppuaiXqPlKiBsWHlmqTgUB8FnhBe7mM
kFq1zezqUIAflT+m33WmUalXKUHOqtdd0635eqO5k5eHI0wiUneaFAdCPFejIHyNFPCTvUsYCHSX
283+wbe1rbMZ+2ed6HIEA+kaaIKAxO0MLoXJGZKiTILw/G39+wS8OT5Xp5tAk5o2LnWbCSE+bBS2
gJ+5EK2PMHiPWhrKT6aXZzTlM7gHQn2cd7Jclduq5q3iY0AL5/AuDwITwSYQH0twu9KT9ez8D6tY
OTgXHwVBQVIcjZSk0pDezZfH41cqEAfu46BpbIxWq3h56AqwZ8x3EgOHLpvpSxxklNmRWyP2EywL
hh6m5Sfl84TE2Tr/AszoeaNR7okijFln5rsOGxKv+24JvMmMM0FSuhl2aSQBSIJPANY92jF+/+8b
d9vF8of5V+KIeaU7PAGqfuxhBlqWBQ4zcc1OvV3kUs3LxT1uBKtT3swa3Xja3JwFUolzJE/zx8cR
z7XR5sT319n6K4xUvhD2naLGMsQ5G4hHNsfQp2+wcSNfTtMsTxqiFGOaH+BX37mM5gnvUr51P0yb
yc/SNgXBvuBEoSNyNyGjUIFjxoLXekSooos7+DdzGJ8n/4NBrK693UFRjkeGOx3JDi5QqThVH8Kh
mJ3tELLl6f3MBhJcaaBUo9AHuCJyTtyLiS+i591GJajt24K1tilzt1/1PoF81irDg54UhB+6aJCG
fO4wGlJXfPVoFFbzGTjI4OU4gKQs0iLD7wQZ3GztTYB+E5MqY/ghXYQ3+u1AOPqv8e6cuGJI7m22
Qc+heGoOMGV1AIgCZFnNAOdnEXSoeS/QxnKGDaA8btg9SltrG/kVfInMjJkd3UvFpybzM8j9zs4i
gLSkVtdoByly+OKTzHRRPrDSoMtAVJ0JmXVgqkVqJjfy6DfDj5HrwLQQx9h5Kdfam4Va8FNYeMij
spsIKGWJ6RcKHZ40nDA+EXXhyD11fTbRhtOc0ui4+7EjzPQhuU/cMKeMSm7e+OFJ8LImQw+/Ufq8
qJL2dqTLUpgM7/BGpPcVIzj75dPF+fA9CELZ8hPE5l8i1ODEWil+6/rgkf7qIzUVCHt43ftXHjD1
F3Yns4n7pkm+hJ5xnBas7RRxixizD9P3kSWO5gTMuvlm4M/VjAtKqiQZQYjkFkTg+FG7I5rlSaIV
4Vj8GyaMp5l9TFTY1Bhl+pyN5PVzhqPDCh3Wd+SGQdgoGy9UKVGKnpGpt5978QaO6osIJpaAZ1Y9
h1qeOJ0WdB0RRjEEzTGaG1Wt1r9Rbzq3v9hMR4ILVkNqw4q+6krIiwTFgZvzRGjDf38b20MTirr3
R+dmuIMn9lgkadbWSBfV4mgsAUTCdbENmy1X1EMJLx9EqhCQkuCmCvZ89lAwfaDTIDmIc6oX/4Nl
UMAntgNyIF0s0IbrVO8xTbl4fSUohEGvrjpiUwcjgj1089urUr7Y0sCmZslzqBHwnKj8UQHp1PvQ
0D4AeMvJuSPOLCcI9r3UnwChSJ+JiiwfHwZLrlH1/hWe83+elsvPMuQp6Usw4HuRkAgKV+X2Peo/
p0N3EQaYbeTKu6usXYwNjwYFVExOeEFEglkhmFT39ArB4zweh3IhzbVfH5hVG57JUv1IlVHgqJ1i
GILU6iNao8AJRzB3Rdjh0MzFVsRaIPGwZ/P+pJMAaLFnxYVthpP9RgEl3/zIdDsyl5v1iWta6brM
sciKYIDuLPBH/hEI3RFwjFSZBV+5vW3PgPDY9DBZjH/FkWm0FDxWfsgUiaUdEMB/mk5113EjRgua
dD+8erOdgkK5E0zKrSO3c2qW9THrbhqL9LDQLLwzki8sWQY8IBvqvfU5ZK3VuJatFwFJamv50lEg
A/5tOM4vLCVq7Uioy1VjGNVG74uyMDU6vplCtNvj6r/9tLliEoD03dpoyeGp4URJoP+D38c/k3Lf
TgquqC/Vv4+3uugECDUb2oqUN3WoG8YEFq2q8xRIpXaSnzFapG8ygKqK/Lzdq16GOi8aJ+AXxlZ0
yHtHBBVt0t26tfGB3tz81kFRL5r1lpIEDsa37FHzOU0x+TMoZE+9EfEaQ74IYmcB22cF/AxD2ACV
W5LqvppKhDWzBDfOAjIY9vi/p+3rNRdq8BnfuP+33O2bQ1ZOa9FMmfoV95DmsnzjNyXrAvmdLBMe
DjZTBuW+ZWPZdqbug7zqveCmyamASgjP/uEiPmiUjHvyU+JYh5rXqwHDYglUNfalNetTq7uIIDF9
dTMW31JA/nwGhRKIUlyObCSkZA5Hbtt6JxHnWzlMicupJgDjhJcYkGrXBzp/q9UuUtipD0gy1lU5
fHGPXdYjvqb6pw8fC2P+btN/2hcGNPYIC3hXxjv9uCtc6pascsnaD7ReJtQAUf04/rm/LbduO98q
/1LahAyj9nU+XLVQqxb3LXXuNKd5RRYJeywkgFzGdW6tz4gnKW+nQXb9psCOjy0cdqksFzTaLlll
cWp70nvacdUrajQOC4TII/0uJLkXxw+/RCd658xcNfWto6XHj0+nneom0jctQz2u2h0hwl7Q6deB
RF8CaA5/AejIRr4GXLfi4t/QDytsL+BStSvGMRrR6NVcv5ZVmsGaKL+4zvWAARHlrYLOwCOq26fN
i69a2QaRDX7+B3sO3vKvgqhJGpJYUswEJ3bkUf9eV3+4Uz/MDCITcWWT+Aue5m7pro1yVEZuowy6
oPYci+uSkoTkkfc0GbB1gpPtPdxZa9/8ZcVoD5EjiJksevEj3ljpRzZocUGy0tRmv2Ma+vE6kGJ1
VFShEYZgunoDqQai7UscMjYC1Hb43C60TEbk5ZZUfIu5eg5X5ooP0yqlPFaolIQebGCUZasKcr+E
vvUmn47vqDHNp3lQpX4JEI83cNBXvqbUaE8FML1ViRmAB288KSdwV6ceZpGemaI6DgoWpdoQi8BR
yGaZ2Qotl2Zmsm6gjKoJl/3F3Yyr18YLgXqGPCzscyOymHagNzI3VPGnD3FsTX3L2kvnAl+erOkO
nr/YQ2SALeDW8VXOY+Dl3GjLhFx14pqKbN5qJP7fB1MAcu9gqAfV14hW2meWd/BALuN6oKgG8m2t
ZWKmskAiOvRhhzFZIth+Ul0x64f1uBI+mqLLtEIBZKgeK+J+KhZvSdMGqp38gmjiZxFy04VSZ/Ay
i3SaLxOidCekqprGBX3mFHXIDLXbxux64800xjOtpudRrPldX2kRJMEltARDAT97/tscRspyf+7H
EqbP69t5O2xZg5oynizgZSaCa3adVwsdEbyXW4B3mSGZb6uxUF66Y3t5CHkeLeZkQDkjxtqPi42v
TGVv7m7YNEwpuoIed8y0426YNUBD5w2+ucLY+BfsuVsZ+QBZpFc83x3cOr1HMApvV7QliUZprkgM
4spyKML7D8s6BX78VH2qWXQ/IUgqhKnkwgRStoda9xyEIgj3n5x4mUz0yfpYJazHidIWtOobEjDC
KUnhOcd/ucN+uoEsuVfvc1jb4AvajYjQQ4QsLysllXPJPP26mkZvF/lMhDa6w+Vs+pk25xn44GzK
RGglQGmb/+m1CGdEdWAnC0icqcMHIR3nVo7aat0GZh4nb1aq39nnb2KfrqHLmGmxKAlC7etO0LRF
cm5WDDRpXw8FHiYxmZagVX9A3EO1EdgaRVQh5h2QuaQtuWclfRK/OxMtuzR5tLXOvm4jvr1TY134
vXuy2g3wnG2TqciYfh53eQBKY6GSp2mFU7IKos33rQXuWjxeAt4IY8wMNr/TDB+aeVFZPozQmhCD
z/LgB7WazjX9vBLwA4fd1OfHN3l+X5H1mpeKAQCHQViQXRxDY92mvDW+PXowzjZaVMh+ydlAkanA
za5KxfBFhfzX4zFU1OALZGItIjr7VC0PyUrlHCDSypRH7kHR3Ec7ErHeQt2/+jJu69tkDL2gQ584
pzuTVE+W7RdcmM63Kd96balnr9sztt4Oe8AvbeYO/6246ovPwZED2tBHtIkTM/cRGwwXxjFWfpBX
XdNUNhkVcubSUohR3EoeNh5sTOmkIRgogaTh+nZpxPQoDxQssnScNpbvipJzGBm4eAarVGGMKvw7
t+P/ycBxZt4v/vhX3b/nQiDhl+K8pXYNh5x1f1MLXdISorM+O7LfBjUPlhxVC6M1K68P02HrVdWr
ND3nGI1AQlgNhfFAblfI7Euev9KvpyGE/sJ6zQ/eYuJroE1vX3TnjpQOZHxkyRlEBSD/nwDBHtdN
j5MPNBO+GaMEZRXSeVcZ4E+aGs72EbkapxEmKfRAgBj++aKxbSLQ/9F4kvyRUjK8hiE8kbjIkurZ
P1IM7qpl3I5VoKZ7gWmvgEXzvtDSgn3rrjT8BObz+7NqKGngJeCHDsFLzRspPGSbAUxEC61QoduS
py86wBkvMWbEy9dPiFbjC4g6sCa0B6Sm+M+jAnLf76QRWHlwPHVCkB0HelhkGP/1n7Nyi+UEWNLJ
cU/VA6HIXRucgSuPcYM9of8RKilyEGI7HJP088/D4kICw46cqJuXR2BFLnoSZuaDj9/v17CJyMMW
KJX2+ondE5jYmjdJLL16hw8lVeA4Ow3CR+xRixi9R1mTay4d0e75K/JxYkHf/hV+wgIfWRbFPAXD
0EknLlp/R+r0Aap6SfUYtncOyRif0GTB1Z/YgSgwpK5Wk/f3xD3h7AsUjLOF6T5mrcXLL8RlcjtA
t+l6eYcLdWXjYrJalrsWXLRV+9darH00A47rq8OLf5rSkxMrVO0mSVyLncQ/IOZglGgctkr8S1h6
ZvQby5ApRg/3ugWOl2kebw3J1juBYjUueX/7LJEVm7bzO4H3AhmZNC2+bF1nVFNCIctN05P7NQSX
wk0CbZfbCqf8Rxn2AJAHowC6nrgKIPB+jQEnVrwVWV05w8RyvFULgTUb+yArXHfRRXkcRwO4m8v7
1xLWZYyXpNlE/pokHUyf6x061fxQjonZeF7xW5urjG1kIE8ciET+egf7xR6rFXL4TFZFnC6FsU8v
tNZsZ4JkvfrL9ie1ZqSF9aakMHkh0jPD/U1zZzRQ+BgSYxUIQTwDA8xXVbv5N3/tzVLfONyd7sHR
pcjBdSb2XIUjQ4NZXPOpsyhUzcoYOiuoDwYxEcySBcCITrXzIYKpHmsc/+xIC3w5z2Whi4NJZrh6
9KihIl/Dm0QN3KDhYSEADsK2spxb7bAs/BaHU88MYGp75Pe+2Hur2w3EoG2wWvJhK6nue7fY5irJ
rbwwES5Qjiv3RTx2ziYAZWDUyhdSX/sZH86chYi2JsXZcHxfWg9Ht2hqTasIhWQnJFv8+qeyxUcQ
g3gbt8X66FhanCzxuxUwp3+FJxRC/q7uNlM/qZRtPjcv6KsfiS43xdnXdC+eXocvCiFoVOGF5R3k
oj4GXSQO995Wpmphpr4fWeWCWp13MFW9OjXFZSsO+Of7jD7ngl7srzt4RUAS1kxiJIB82QMnzYAU
LqjXwL5BgE5sybHSBrzGxPbAyveegU7zhEykv21+2u4nQcTBpeWfHGbPyzVrXUKzvDlstc4auOx7
yTLv/z6bh3mAl9HVig8/XajmbquO9l+aeTGT1eLEu5BmLWy4SKX1qNTTSkBfjvKaDHTJPETxDQD/
0l5s8qslkfIv84INK5gL4GZXEmtGwTkNMSmyVl8s97vGWzVU6THgzsRrqQOF0iB/OlYMZaKXCt45
D8Tl0Gohpdu3BIPoMrE+Yy/cDjf14sykRdFH9sPXFP40aca9wLunLePb/BHxL2bWKPjWcfmECPmE
j/PpOjnXXMLJpncB+aivT2fBu1atIgXt5KuJS9vKoctE00AH6N9z4OwYF61PmgK2u4cDPwp4gHLP
M/ksUamd2+WmnbhXEm1/ieOMX5rEGbUYrOyDeA84KB0kuhSVGNpjMXwrQn+g2kvgQ1XWbB9eOFly
19roHnvMGjLL4TGK4HZttTVfFz20YZyiEjALAWaryNzpaE4+cg9GzB8NCrF1tDEEz6nqkdoqVsGs
vpi2pJ8MpntKRbojxtySVoi+d9abQERcudevu3KYdpqGa1KCDssHDDZy3WORSIkPHF5kNyYeQNX/
nup+qQVNz/cUPZxZrgC3Nb5OEZLn2vjZreBxj2nAdE0KHBTnOdoZPnC8T6n9Z8/BP5gs1HA4Dv0M
GW4cDjZGPRoIB4G/tuJaZTDoGroFNJIHgvvBNKjo3qjhzi6TcUcrZ/3IrGeYNr7V1VJiJx/+lLiL
+R/vnTEGCpu6Yt6AcDz8AS9ZhQ6GEsgYmV9RK6sXjeMdwQKS0JY0PPLubtattemkgEZ/v+Z4FoFy
9FhmykZwXoLyt9n9lYnDV/cPsHZuS8jI5MGd+CnvGoAlp6mupk2JHoX2qtv7hCStYxlh+efpP7Kn
St5pF9Bx9UD7SWmyQsTGZNWDvOyGrfL+XLu7RjRECovpfOBYSXpYc7zA5jS0/mht8qZEUHTFTCvJ
9pSXGhiT7ASjsO39yKHRUB0pIDCkvVcngcDN5Ifx3z3H/Kl+bG1HVRgVmxHHx5vte5PJq/VwtEYL
UN+VApzWEmIl6Ar3G/GiSqdbBYPLlDbOzHDki4wehvmGGzfZhgDw90RI9Q3Ux1AXhP28XoJiJkbc
cpfv6lXyuPPh37YhNq6K3rbegog5u3+kipirty/hRI9BU3Q4uKd3dyp8Z2Wtj25ngfAfWmfSxTRV
hezRIcm5jCLnzFXKviRDFxpyx1Zn1ZS/xvIP4W1ExcbdrChF7I1CEzuveW+Ygm3dF/aHcGhQQfMl
WwugJwPC8Yw/ntm0bkxc85bG5Qp2wjcTstbMfvtadXDedU25ofBMgL+3sX13aiRLXCZoWjqS/50F
YmTdpFBd3rPquYqTWsGPtfJxtiLxyCzUwJxbqJW3epNqNBqsm5nXHG92D3rRpP2Zw0PiAJW4qv2K
Jvvs/HsEUrvgeB+mSbhRkr0+jXckZumWPx0QyCtI0BAEdRpVcRUdU3Z/ytValz5c66PGcgJi9Z+A
lmQTsMQBeqc7NGug1D3WNm1c8eHm4FAbCHHhAExQxPKXGY3IR4/ps7mU8V1qVZ+WPkj1F8kgF+ql
dEghYGwyTZGNg55gr7O6KttByF4ORi6HdFkH5PqCMFfOhKkl/Y0XNQXNIPx9MoHl4RcjxR54X5Fm
VQaOW7gppisTZ6ozmNb3xh2QO5RmdLjLpj9TY5BgdHgyth6Gli0eWqHgZlFvfYqSDymoWzcFSBJw
pcx1E7GkzGYJBHBwApSLv5cYCL3RmjiKE5oDww/IVkFvalcrG+C1exYIZAM8HRg8yd+MdqJFIT41
DTP/xHixj09zhkCQGctks0TjVv3Fu1C5SaEYq92XfjH/0LoOgewWuupCQFgzVUrK4titCRdgMhnh
zv9zvt/COndLa5z2rpN/dTmopIK0ecKp/YkTvTbuB1ryVTsLuZUXjGGRGD7JZV2eUIfB5mbhgPxO
xnuMvGoBspkWYe4pv5KCzb3ANFriVeKXoGpAEjj/usSmcaa3Plwh0i0W3hFrivjrWv5qqUesRouV
5G7FjVi5j7juS73Lqr/RGo7DVIhkMLeUfbe9DSE35A5l0lDzHz3gmIMsIfAkWN0PbsA0lGyvG74C
dkMQGXvWRrMtM7qiOIandEItTNffo3CF5HTEt+bNPlG25N4YeF2aziJaOkl0NXJKXMDAHVMA9xye
zwCJW3mOoRzaGOl5ULIf7Arm22QCdqbLmGNJCb9OFwtzJN7egpj7g2ESPLZzE/NVYr36UEwTwtSP
q5InfIGHnSZMuNO9TPWbyTIYu4oZEzFrq7o9n65ryeKDhih6ZxiSMTNHfGoAuK2SEhL2uac3KLGT
X9X3fq/rdjPYc7NDGxMjV1NI86gjAoVw6w6ZWSUM0sVqiN4srqLSe7AcgksQhX77EvHChZq9DQ8t
uI0Ww/KuGS+L03arZtGeIfnBWEUOPoHtIx76pOW+BBOeX3PNnJxRDLnl0sLPViMmksQHMGocgD77
p/Wpwtem99+vi1dF9C3mj1+69GyWQ6Vm6OQQ46VOui4iapYiGXbujlaSFawOMqLTPyKnNuigfUyR
lGBg9uXTSimKvvxEdWOOsZUD5QSeQoc6svG9rVCwSVisfXMZKBQv4VbFJcCuh69CBl0jXRJPiVTu
9T3cPkAUiL7N4497ZsRVwKihVbh2NDGGe+3Ryuu31n4OnXPFJs0ZIdVak8HA9Toz+YVNfpnne39B
/1EB8xua3/+TCJiVldUYJWimDwAQ+qoYlF//1SwN8JvlgCLQ4EfwWOdMeOECND6BHW5wm5fzDsdO
xXUzZUHQ1tsh8kDG7S9KI/RgG3T0hKZ17H+ljDVxLoItX4P7PFnmqs8gWDwMddXFHoqD/LAmQFxH
owNZLgZ3CyLJ3yCA9J6Q17J6EFGkaSum9dfOo6OVED3BER4XvAByKGDMaLhDVee0dXBGBy4CImKs
EWVDM5hDoJ830zBAHUtBk4Vu2QBTvYcFn6fdL6HG3XVkocN8okJ+1N83zDeYoHPf9bMERJUbZ/Q0
6g13OlfFqkBx4b+LMnW3/Lbo0k7j+1LQlGLr73nKmSKmiWTGHI/aW3A21+xbOuNrbuoTrZB7Rt2v
EgthDXEJ/n7v7GoeF4980saq9NaYcbcYzo8V/44aka4gYFVXwlcvH/5v8KMpsAXraIfoaPidQVh2
iP6UmWkz6LQTdvBJFnPLROiuVvz1bpjOutvZTai0DVpT4ljSwxRf8L7v32PZUYPTI+o+6oYf/CdJ
sRuaQbrQs2v68fZvo5k0o1JmG76UXLbDXc/xY+jvni5ahBq+26VdA6wr5zkKxtuOZPTefZTaoDa/
4OzJ1uQ4kYFRgoVR15UKF+DUOlw1d+Vz9894IQh30jY4wG/xOSm7ym9s8QacoPV9idyU8QakXwLj
dhNVKps7w+1WiOnu4vvwB7ZeY7g7HS542UfUO9+A0Bu/X4Yy3vZtaZuMqjBSOi36SZ3yTybuG+2x
4iwy/ueg9QgKt6eZVyeXbUTKBdV3dLruE+oXAz3KLhK4TrxgIyGRb/TN8JBTu1drz0oekZeaVWd4
FWUUGlu7PxqYy8QmQNEVAn1YIk6gYvx6gU6l23WSQjt5/s4yjWuZhrYymM+FhxOL/BqYwnsT4teb
BVABalQ12ES69qd7BRFYMN3Lf2YLQ7kRq0eRu7844q2ditZccarXiJo4BzCrOBhYc8Nesl5jgSQc
i8SSm7c+RCzL1omaA/m2tGvmEXWv7SSIASCHsa4yhhQvbLl5T/LTGTkTglEk7ZOZoceJLQxWIOQd
no4q6Y+OlqSpqfIJr5LCvHQmBReTL67Q31/WVuCcJWmdqOiykuXrDnmJFsWkQ+OVt1wDTlMacMfJ
bTYkcDpcYYf570I3zO5wUh10lspcGOcRWHq7IEJxiNUuUPgGGFliS7+NFfWXV/OGfiVcI5sscO+Q
i3QnSKNgiMBzFsefdQJadhFKbn3MZV0IADHPdkn6fBECd6e9Fp8u6OzNMWiAqo5PsaYsrfqHpr0R
2fXMgylCA+6SHn025WzGWJrD8V4OsxemOoSdHw4nposc8Na+TERoAopdpQmaJt6JZWb8Dk+P4Vzs
0uUPMyFbWLTmxRekMx1PyMv0It0J7xk7V1ExnhImRjkDDbyks3QrS7rFTzLWYmqkEjTdwAnKJcu2
TzKmHJK+Wyw/dlIssuBXVsWhIUFV0A+a88LKFH+vyANnKl/p8OAbrWCWWQSHnWlpwbdmFG2zcHA3
sXsFafKQiitEa+LCQG4aOHYzgQrwY1/V64Z3TiGIaIDYS81+q9O4armLPZQXpgEtMdbpDP+GwUHK
6WkMfHJhyzVFNvcTJ+nqQ/0LXmyHXi8tDyoFrIIGjYkfwroU12gbzjROeqoKitxhgEbrAEgUHHXN
f+Vnlixg8sZ6qikV/Vnem8/0bjQWBtptltjzUbk/QCNawwxMqW0GmQqbc2xBEOub6ze68TthsD9A
95UedILNqkTSPlQS5SssGPLmDrFRVW6V0lrFavrwx9d92dT9pJS0yt9EXjsKLrku57JgVPjclYao
UfvRtv+3uimfKA3912sdGPYCuLY4dJRqGJETsp69/YLV+gz/wqDuxhEut+AZMyJq8mOv2Ag8t2j8
HVbxwckOAz9tCC8e/tLGix6JAdwxSQgAfLbVcqp/KsI13M7Oz2FL2biKmDiFATSJ/8PvfgIgOJNJ
CLDu8D8fdrQ9XgYLHkUoaCkGO2/Gv9QM76cpwUOixiVONH1pwM3eq3+HbZO3A6PKDN+Wf+FBM+46
KI+/3my5wwAeAwrw5TMPJrpsw+KVWPPnuglF9EtvyzpGsv/5I586gI76z8Nc0MK2O1Qzgk8RZnhe
/+DNAguneKhgrJvAvlB+TNrBSaE0D2TLTYJZ8JO88nMbtDvLi1nSnvQ9ZmSWTerGyx1vkYYx/iXK
cQOP1gw+1YDo19GsqZvC7WLC5LrChL0SwgEqEiKqnRkHXRYH9Cu+yoJtCTP7Q+IGae8pkjSIlEO2
wml5oYI3Py+c875LWwTh4WuKRzubIMrrMKbuNvmknVbJOfE4nBF23AnrKEZdmQJ2DMHuzSHrA+Sa
U8fNqG6iBisv5JFVfyRfN+axTcNe7QTpHVRtL+rLA896aoVQKM116oSjQCRwbv6U8tUWznR2G6eR
rGqeaFhko21nAyHjkq7pQMJCivYdGsgh6P/Kz6+HhJtG+6453YgSwi96EZiGm44LQ0Ue2GDXZngc
V1HLyljiyQWGS1xT919s47i3+RO4SNIFmjSHZ9wfjFdBxnndOocv9DEnxj7kK0yiaUhma0Id2feS
7akI4F/6WENE0XnerIgVUdecSdKiFQ6zZJKj0KXb/GPxpi3LEKG79h+yK9K4NdPXGVHMVw2xwdRM
7Z2f0+JaaKzY4Zh59MD64UkRnArxJOwV+9mWFCPqS05qWU12E4CBdpVTJUVhMyrb8jvPwFIX64gN
7uhpomt5Ptrkufw+r4Ds5KFJaDUYMFKjb23tnvYWPla6RvMZ7aYKmG5AshYCVf7BpH+7yqMxdUvq
NrmdzY/lZTFGUf1ylmmawQHBy7B1VYWwOkXMz27kGJibMl/cw3vNqVAjKf3XLOJBoBxvrCb/jyab
bkzuzuqraPUZSDh76J/8xIk7aVfdBhzT1Ff5Zptg/UdxEkt+pxHo3P77pExWzi2mrl5jsZL8rVFy
hyJXZjhihlmsUS3TP4B8zWQOAAiyl7wZt5cGPOMbrO+TPQ/u0T8y66sT+tkIbkmEXztDVWZaWniQ
QKFByVB7+nQM91bmlWDXV3V+DuSlKTnUMC/8bYY5AYnbnQXw2pntopKlUazb6+Dgj/1acOZFvokk
/XlkIlfVklNc9F8sZcxw00nBuczTRhCEHvnt0WubfSq/pd3cTDAduGEKzMYALTMMDUiZfIRetAhP
BFNv7/IxbNV0tHEIiX0Sd5g926l2UtdseUj0b7glowOXfxOD5KVoNsoc6Yu8wJQPUXpuaSQbA1q2
j9tzsnOgeQ4AfsN9Pu+OX2cubhuP+bDkzsXy/8ysvKLLMH8oifhhmjbZ4aNT+SXu3Cznos+1Hwga
8D2jCXfd3NZuVuPxWyl5MtRfb/MXyrLEkQ0h4SEv0wAjpJ9QBivabhWKJWoQpQQpCMgOxyzqYoq/
AYCV+ZURHboNuk+BjOnn2Jfi3N3gkISk3NBIBC+tfS/U3ZPyEJLNxRG1zTWxC46tMlFcTNHnyumT
EvxFtcHcqb+rwDP5bXlRtt/woMhZuwbcvof7AXGuRPgQrYADUxXf0qZ51rNFhGm61xNZiGpUzw9m
oYs9QsGW52UoGIf8QiuUIkMTSd8WDF7eua/LdctYIY50iMjOXyyNCwYiR8TvT514a/PzbZfX+VLr
GI9Jfu8TLHZ7TMum3kRMVkiZ4Y0ehv4YZfRUZJ9yc8+MSrNemWnpeyKHOGgBsyRwy2iDBGJ9KxlJ
TNO4zdrz8Z5J1LYC/OGaHUzL/D7FlHIm/9amiaaBTjEYwYiglXCTzNVanMUwRD6CP2zJE8sqdds7
MSkrgom1v+UhWTvC3FxbK28O45KI7tUgKJ8TK4vV0lmQhbT5dIeyEzwhZz1N8v/EA9sgSovwGaCe
Z7CHSXUjW8qAhdg+YS3B9X9bg4IYLP4pkY8JIoNnS8nkN4MrXegaMlFnHMAnMSf7uADSJqGEVDG/
5BLQTrzFrfM1zSP0O/iBlz/lUtxx1UFJStSnS+nUFwS4YQpxgKSDb3kvQiIOjhHfFeX6GgQ/NdpL
wWQUvz/dYfSj0ODRIJHq2p72CDqvW3uGRRMaLM/pMh4Ya8jNBeJMnG9yO/Cf/cc09iBN+E6fv7QL
8qmLWkuozaeJlHV755d04QneaNwR6+tUSLmh4Ni7yrxM4B8KzyrVXyQCuu4eF033QpGrnAdutYI1
vD0jJNXe/NrjDS8HV3saHOSSU1OpagXZp9807fp9XDW75l8xJH8RRUGJZorZNWkQ1tKe0393kqg+
agJs7QB3/oihnjypNKvmK8dNvu9t/zaE7QzdnD4aBmRhIZpt+E/PuKNp/EJsKTgAj7+3arsFDd+2
KgeCQG9E1VtL+dw9yYjfmywbfk6sDna77NU9xNuRd2Hd0gJILt70GFJDb9fGzhpN9hAiKAo9UNcj
cWh0iHO9YoeuaSFrZ/iL6wYuzcbgjW6PUbeRSkI5Op7QbgHPvcoi9ouNz42DBqN74YFzu9gG5bAe
lcHYUzH/dRYJ7/iZ6kExm2dh/j9y3VwpxwvVcHLqiWBPnw0jWDAYoCxaBB5kzUa5Wd26uEMwBTjn
WPSE944RjsnqyLi1Pac/6+L/cKJJ1hhvb/12Sysf6nRyTKuJ48slZfKLpRVxNUzVkEBg7iFVXe/Y
UXqfAf63hMNc0tpHK7nuhuwPcVxWMj1RcWKbYyi01ig/AQbNkV257fAgYqEdluAzIVdiKMHFel4Z
TLxtb/JnJAfzOv4rf8R85trI8hprpTPpnU3paD6p6HYsh0XFBcswCFFlJrllHjFnexvO9e0/jFsS
Y5Kq+cW6WVCoyVU6n0g9lQh4REDgv+F568089uh/Sn60C62LwXUF8HeSkiF2OrcuMBji7ICoyp73
Y6l5iPP1w0IcEK7eEL2Bwa5zG/yyXE92zrI8Y17cGHEEuaFcG45LhF+e9ExC2E5SB35F4oNMVSKu
vBryZI1CNJGtmUZUPH7u8EwfaEkHnXxYS0+XEE5X/fXCNBHQG8u13CrjfcR7fUMUTTz4qeT1lImo
RiRSQnQO5bAlOVoHoaZQKrOwwJus+ANgISfX2BSnfqPC0Tn3tC9nuvXPJmJrAugRwjlcRUIY9a7G
U8IPc+1TX7eXvLglbC2NMWvCL8KoC6tlzX5j53uIDA03/z34el4yV5qED2VaUEno2KoPYiyg4oew
Kn6Os9SQcAaCEvBPdJAy0AuEwBLst2gzIBdfdGJ+eguyXuo2PPrPdymaT5blM/ZnAi6UG5f3ICF6
UvGoefnStDVzys4ss5H+gvzzbJzlxIUwOmqmcpVFTdbBnAwBJDeaDWExBarXGZnZgrciT7rT2+hG
OH95T2BhtMmw0lSb+oJ9EnaKhEl6HxTIZAUzPHUrEULNWB9BYtwBlvm/SOjW0BfRNFmmwpCAf1cI
w6Zh2Oxi2Eaqq7z6YLnUrSj9tprj/2XdQy7iVIlDAB/ws1sv70YrrufgSOFDg9qcCzKFG7545m3G
B3u1xajyY4MFJO6D9tKz0/fuBkz+toPolQI5ur6aMDUi/nIXQSKlmmtl+zsm3frkXwwKl4rrUVUn
YMsc+o+xZo5qYKZW7iGoNoYcPL27YMd33AGo/WDa9w6YUoH9PAmJW+ICVcVZyLvcJ8TUGoPhMtE6
Uosomacwt55KUkkCgRfTFMrjXxWzNLOUdLEHER+MGgJiJT5/lZNvfhZh+XDpumWkoIu+D5cuezE/
OiwfjfyiVd1jOBLKq9JxUWn/VNVsybfulPM/PxurXw0zhSZHRBCsH+8STUY7wd0YSwEfpXfxViK+
VjfPoH8fZ21gEoL6zYjENb3LU/s/Uo4W6zl13bVrSJbh8/AVTWOterssrVNyzJz9QXWG4VGtEc5a
Hauya8DXvZxH00vy1cOi99VuGmkkzRb2ODAtQKYFG0isvwp35iZEjUpYZJR4TZ7qv0J+C7/VYFeS
YifOILgELy9Rri7CxE/yMRF1bQ3D7f95bpAGGqr8h3Pj+8YayXvxQWJxTanQ3D+bYBPuBREzqgbV
yXstxi6oc0EIffbl81o68f33YCLaZxTOt0iLoTHE7RlMuLaZGER1GdJYBP0w5SvI4oq5BzvOwfCf
enTSBfVQhFQgDSXB2hVirCIapxeFZUiNAb1Y4TW8AnyD8Dv2iZ4z/iBd1quW3i13gflG76Hw3bga
Cu3o1wckOSDGTS+goZc7eLsd1ZfQ3nF5M8wRooxTKEAezycIfxOo7Z9wr3FGX2aMZIZl1VYSSO/S
j7lyAOHPgHZMB7005gaiPD+NM39myTbkxA/Pv2/ysrHE79HprdlIoE8E31zGlFVw4jsojnFhGolu
uFvBiYN6rHDsQQU7001x0dzq24uu1ZATkTq/Ks6+xHdaDdtWIL+DRlMphGXbbhjx/Csq3ZdteWY0
VOe0YSn0GkAmpO8bR2CE/4iYe876IASrMm9j8rogxplht+39DyTRYHhjKsOVdqT/c8LALbltaO/+
SkjKFHJ7yF5u5coPihM019syzsUJHOqO0LHgAz3+hWLxSZCXXN2E4M4JNxy47lcZkzG7rG4pY8HN
CaKlchyUsTrfylkKadKEqU9dyb1Jkz//2s1qta4Jw0BnD5owlpTT3e7q7nNXnV5i5tyWx0A9zxiz
cQlJ15yMM1iXIFjJUAk5NiEfwaQLDoZjnZavfY9pzoTy2h6V8DwwpYppRfKYwOo9f2E/XNlRlHwe
+Kt5fnNCqAw26spFEqSvL66y+D/5ZGV5NLMpl7+qhHqoej5ZLKOc/+8u9h1o8n1vOXtGphfrmjBU
dpCxB4AwLV90gkfoS19tOE05I7unEi8dbEH0W91v+eKf6XbdL2tmtHiKr8oVVxpMwE/odnST6nKb
BOhJJ1wNwFSsRHUxdRcaHbtr5nQcWUlJfa18ULviaWKMwO5wA3xmswJXYyVHzfmBPynaGqRwWxUP
WXMKYVrCSpNIehI1VqFCCMHXHU1aiV7Bp9cbahgRK5wctUlX8juKFFLSWWguQZM/EstoSqqnfEYo
H/Mlc6o4W5ALrcB39lux4XcvrthooLyVthT2kpt8FWFO3vTNcEtX6uqLv1zyxuy0opRLFjp/5Yuo
yH1lV5wGgpRc9vL63yX/x/qwOYO2/xO6evSSEdDxkZDz8B0R7/y4wjxKea7ZkprCzEay2yr9t2jZ
KPN0XXfcC2q3U2xPCLuRfLTEOuSkKhdX40umWJ8u+AtwSwKjpSz7elv+kEfdLnz/4JlS85fhKA5g
5B/l02vpbJENKOLajUOvo81p5TpXKUo3zCChFNdkPZGrOXug0RPARq/FkfMviCiP1ykUPzBqpB59
diRHB+Ihi1+FrGFhvKefpLpOJIIH9kHvn7wsRwl5igExX/XWjgqeFAxQ9GsKz451iDlr7F13u6hz
6WnqESatb8Z0ACBWgwMdWMjTsfVLmc7HrPbCe3+EVD9jAROIRH3aLTi+g9qp44g/wY83YeeqcSn3
GbUiKxhcV9hJHeXJ2nQGTFjndkHS9BxlIrxtYNN8VJ76JQU9DVaRNmrgW61H6KGcX8cbgBYadHrC
XJUJAvw9Cm/hosDMBxHxxVc9A1t++vDz3J3kxm151acINZ0JHbZcdsIsC8Eh/dpxgwYJk+aP3AS7
5pkjV9HbKnVrsF+AlEYuxgkEpii6EAKti3w6MUC/Ut6HBLSrGVyCkeSIrn0LOlqzOz6XOdNyt8Xw
p6njgQhyGGIBrwpLkf3KMRLhnZXoUYcKIuJ7h67x322G5KjdxB37A9fYAx+29kszRof1N80+AiLY
aw0Ez8Vh21Gym1Bf8GVuFRYnenJ5r8sg7fhFyrRsx+srgskeywZ27iTtSffw+wm/GI8JvQcL2m6x
0BTXsAu7fUAyali6NyA3AjvP9erkKMDYn0Rwt+7Nyf4+d6i3KXc8gOQw+q5gt/nGNB3xLnPo2Nvf
tLphfHKm3nnN02QCQ8Re/z/Oueee6vYLlHuFkEd/BqqukFxg4UkMd0jegPjofIXrKWdvhtYDRvfQ
fJQhqpkjQdpAg7epkYHNoGqhD4Aqnnh4Yv8kGqrRaHX6bc03By2COwfMrO5hrUFbMBZEZeXgR700
Td8tXbO53Ql7WgX0QrH9B/4FB/2cx4NWF/Q0KxQ1rkSFticG/YgtcChcLob7H8nBl2Ypd+jXLdEe
1zPg0tOYmrNez2AlwUvSHO2TpLZCHQR1dHNxSOYDFvEyB3PIPfMLfjxGh/xU02flskPwX1rPJuEB
3/vSrO9II8RzGVNMhd3JLMvb3Ioz0SKE3i40YsFnRw0Cv8SyA4PdyfTs64s6llFW2ufrrc0OvQPm
QePCuY9I8aA6cy78ZTnRRau9/PBlKKMIlgO3HK+vDPKYwsEWplsiG/nMCbwNsMMF0FdB+7B+tRbS
I+QFABZhQaYV+m/oPK6fOnmWOpweKXHfRqyuP1IyEF9FUN3UcfgmOgfqLDcfTKuoh9mjpZrjC9KB
owaqNINFIOD5TZzh7DCJ1UG1oegK0OS769cIyelMKXzBqQWWCyxhW2m+KNzGdsDRxT3EbDfmK5Fv
lgkwqNi1ZC/mFD8nrlZdK3TfbQLH2OYLfj0sjuIZp18KDNu8QX1zL0VEHOu0B8nXJaRe0n834jtS
8bv07opEc+IQ8WQCnMUWrXWTexryB+jlNJhtlxZu9JUoZeqIzAuCBKIUWjwmg1HAgZ/c6EHNuviN
54jPLq/MrqXWpOcxyvTGcEilEQHcX0+qC8u7I1NjWi0Hb0F3ZHkPxS7LlBJ2j+p/ylirWIsJucCr
9W/dnojU1b6jEXUeXRaKofHzO1IUCi1iOXiGi3xkFUy+ePSqugw8AE7pCBlAJN4IIZ7fFjRilZ77
xyWgjMEYxiblZr8NpmXtqE5MLHJqhms9h9H7k7m47xHcQjDn2EnAZ1sENhe/W9WwF6krtCg2fxcb
8Rat4NG06UpBlHwssYbVa5WiDwNYtlGU3uySDLy1Vt2RVr7wStyj2J9bOr4/4BRHWCS3URh/Z3xe
r/qFWbkQyp7IMMv88dQz4q6xuPwKio/F/HAQ/T23k5ZfN8fqQNt17nCgFsoh08pOAm321btNad9g
4ElDkLan8s53kRLXMnfEperqLYgYzdHWRI6TC1yts8TZ0zbzW/Ttmds2jfErCGU89uX7Mcs3koLj
lhF3oOe3EZdM0fjKjps4wL07a1VoyeerpEWSAnzOx0eRFkwfnontWF6TC0ZNRHzsBrDEtOBsWq32
0j5rLtbaqUeVjwCNlGdhtzOiUiezO2kD5VgbBFWwLSYg1qbOYAIPpxiSDUOkzcRLy4emrxTbTwtG
P4medTa7J3nhBvk4y5X5BtaclXwMk6est1zrWcJGIceGqpTx9Phv7O/C8PgnBEkZ1y/JKijFbv6E
17TlAWQWYzRc46E1x6634fwWX0sGzUhI9rRs5NrgjItXAH/RZzvlMn5gQR8NlOQFBNOGcQcBH+Jn
jofZpiIpnR/yurw/M7dezYIMiQnXd02TShkmi6OWj5+USa8su5o+DzQTP18O+yii4lbXLUezulvY
98AVdN4AnaCqsEv8ti7kIziobEQyEXYT4mUIOHC/HfE4+qNXw7sPDMeVUmoW5QPBAmeayMNxQkmX
iF/OB4QQ1ydLW+ATU9dEMgP2iKUtGFQQU9MC5GcuS/6OytDyHimAU+AcUhYI57vh1PpJMZMzL5GL
xYA0zvqeF30EB/r5oGalELcymCM/TO3nIagKm9E9u8w8JvLIwLf/dsIna8fS3ZWq0I72MWMxNVNB
Xbu9SpTxzk2U1KSTn6g6pFdvAWeiRcfVbUtR+E49Wjr3Ep5wOO5stdXqEGAGjkRJw1H59GloLCvP
M3wrPg6I6WHZQT8MS1sTnp9iq9o6Klg/jA+ZRC9EKSOufCTK1BJkP2toHLm4r1kfigPyydNmQNHm
A7svWCLb/Hqz77K+MAOCz8Y7apUxct+8Vlf8AkX2gwV/AH77oedf0+veZHTkWUfoSVfvbyMrbHyv
Wsh63/Z0+DYPVkchwHUs1FkKQjSxFTl1V6o3wbWvNXBCG4VwD6K54G/DIaGAs1ywMVu/6NuShp9B
nSkJD5i7eTYTguezGRGG8LwfJNeAfw9Euf0FjeI9W+OdIuml2XNQBm/hYK2hyqf4eeePvBZyXw+Q
boiz8D9Ypg/+QUFmNRsJ9IZQMMmHmRyKi1/NWU8VZ0xIWqc0Xe5WrlHO41c4PxKpswUfXCKNG8zj
hTgEXImKmOJNNyLaPTnGYpGWX0TfMFlht2JhHF+SzshUZK2PnsriMdTCs/qsxPqz6sQkIsEZTWKv
kLFiRZ53XgC9C+nXzJrbV8s57XvQ+nDYCK0eLa6dOhiqjzLssxmJX0ehu2wioWsxjvcbvTxW6h2E
21PwnIpa/Vm974IpsADIAuTZrt65G439sJFPeRSPVvJvfQwtP0FACIrkm66l+9wxzdH/Ez9MdYm0
Dn2gY15bVa0emmkEufZzD/yeIuRWTmTeNOvfFN0jtZJ3aQaCZhfuOjM8Zz5hEdKgoiJc6eDdMAyQ
PkHpgPylorV4j/i/MVrL6h696imnuJ8HseCPSwIVJNEJxI43ntpLZccT/WF+47S2rmlrN1MluPdB
qZrv997wBFb+86JyW194Q842I621Bf/fALGTUUxk6F6rJ7mMr8SQIP0B/ZMpy5vwp1tTojQIBwLE
o6W1GITaRj39Iou30mV0GCZy6VYC4z7NBQc8hgzyQsdJULTfnmGviVLt213zWSNjvrPZicOempF4
Wp7mExMn9IEaH42nVWYvUxkKCFkE3y163NFvmLdut7pDy0LydZVVCCPC++BjHBxpAmG7jPANv7Fq
q1gH7NTIdxNNwz36SRZefxYwUy58A/IThngZ560bj8diiwSNcrGxBMrAQbp1FHHU/TUvb8cMPhRs
AY+dzwvB1E3lXa07Wef6CfCKkNzvgvtffJ0rMNRUnK+NDVz9QuW7CMLOL6tLntX/KyQqufhngspD
XUKRaqFbY4Jge0/PLht7gMAiTrlN1LUoLZfvTFhRPS+9lr8toAajUbugiieefKQpmQJWeTDaLeSO
NGDCx0xhrqTFpJJSH87wQiZ9Fi9S9KOwobEpLD68kNJ8q063aTH7PXW+vivjfAkr7i0++WVxe/6O
bympkyPC7pajriaQicTbyQNtDjflaV9w+wdMGH5If6juTDphDdkvvctzNhT/OfsFpqIlXK5rN77n
CZTINf5u05Z8lZ4a6HCz5gEa1VZE0FhzTvhv0LpmUdUT+JitIm6uRAv5cPa2h88F5kNCdYvHJIUt
AgYoYw7E/F8q+mf0qWeT3lsnc79peQTFfrhTjEpBfoyMPKRE5i95H0Dv+Ek6DW2dUhTtAO/cTrD8
gnhQ+QUnxmqF7zbR7HLt5tdG8FCi9WUkxArCfpKNdTuqHcgCXvrs9XTLLmjwyRPRG+lYYSl+QRFZ
s7tBxeOKEpOceUTp5b+r8FElVkaznBksDS5fMPXqO+D/trLdRSaokyRjhQfEl+4XwPTA21nVHqsa
2Z3uX/O/b4giFkVpwgII5gUWuVkgTgkNYbBaYKmvwU45cKU9q/fJaTgQu8cPGIRCLD2SSSX/STs9
dn62JYBmmmCSkFGLNo3zy6+Rn5f97hhctwmaiKW8BXRwvZ41t2u+yJhrElYH0JDrOT89Lk/syf29
z0cgslQHf7LlQzCXza7SLtfzenv2xPR7ed1N1tOfIoOblAvoK7k1eA/lrTQy/6+38has6vwaLEF0
c0Pj8nzf9yx0hq2PE/V0lnIS8dYH1Q4dxN42wC2YPXHBGXNRTbSxLeZ0lPBxVpx/2a2hrWRNwjo+
b/CzNG4spatN7W6yOZYtfeZ8dPWHW1j5yzbGWtYmw7k/DNFn4kw+fenA+LVA6e+wJdpB+71Jffdo
a4tSgp+3n2RYvJBwikeiFs1t31qkh0+2FRKC8H/5QZbgup9QC9CGui2u3OSuzqjCDRzVYthFkXrw
MJvPts+tb0P2JbaEeEX5f2cDrKp+kWS6X7cwiFduMUBKLmjYdx5kf0al4yHm8Z2QJKWJJOTCpxBT
ZcDsxYuzpcVVldYtEH2Zzoe4vjKfl3DyqCGnrJAsKqwDR8pNXjID4vKrHOKDgqeN/di7bxE/+c2w
GCkTdferRCft4Mp/3SGX9FUXaebdK0IhvTT12kXF+4y1TEyGZOqefe1YEEgba1frUkyyRKSY8FzV
R+I1WGQJNYI+5Y4kc8GHW1fyIDbZoDZ1z/NERylMi3mj7ek1t2acrDHuGNnEkOwyzWEChGWyVCUF
emMHmylW8ucjPb4N8Dh0/J+3pl0CuQOH8+vxYRVKe5dBLSodWPnLu9UTBzXB2pLH3iZ9vj3vEt0x
5+YEAOzJW7uzuE9w+Ku+dSCDEb+BoK/9xFQdoCUzGzQp/k0e+acXnzp/L60aMLNv4fVs2/RUp1Ic
XKvQE9WcWAUFiW33nZ0f8ddu8bEbVkZHuCMmdwHVtBQXtfn4q9HJZzH8Ph448fHezPm5WXjl64pt
g0/ay7ddRVI1+vw54l6bpQNyfFXeUBxdMuIUE3FEA4TkrZp9Ur+NUy+OW4NpLjblcEvALDj5L/tu
KfPkM0mSrHao1NxWB/CL2j02WBpYbdLEcxIkE4gL4JdJm5DDRJQApRumi4g+s2k3+L1wLiw6ipVz
6/Gl2wJx1qGfXVo8k0O7ZBr59HhW+ouvZW5YJhnAt02DdiIAEAkOVDHSKIyXTkfGFyjQhUm9oKGs
AJ0fIWMxlKle8slnCoNpc5lZHPqtzon1I1aQhrL2WjuhwVGDnxK877x4Y7OCjNg2GyT547S++KSw
UwkJijQ8dnlwZjT0h/J6/zN2z9ZDITO5lqZyr5RVoshDkJnABvoccdYU610/T7mAKNHvZ36RJh2+
2EiGqBmByukmMFfOF1J1/bfToe+4ny4Zx+zsKtWww2WCknqMe73YDm85owLZHKXAssDhezmbBm3w
D1PIxlRpgzOP9RQ+BPomNqj+YPoljOkPp+QkQvfVd5jXR8lqrZ1GonmmyzxxkflueaNDWbByKyF6
CYh+yMJ7SlbxEqLtyn2UjPvhqFcdTuurWUWeN963vSAdJy8igd8bmMpK/IoGHkHMmqochIj6y1Pm
CZSDkB+AaZJqH5oGGREI6ytZs3Kp/9At8jJVzG8w4LrrY5ZUXNcna/rWXJ06uTdxx7r57SdUsghA
Q78w7RFs5xCj4Jcd21Hb6x97dk9M9ssMqqHHVf+XUcqa54+/bbTzrlZGuQHSl1lCduJOAZb/VoMD
4MaEX4MnwYgSHEEKPn9JGNCvcHVz8CVJnNMKo9ixLV0snGSAAm+Xr7ZSyW2C1nzm820lScOnhu1U
lZeOhkTwxehqQyj9bEi0EsvnGKQH0MdEST96uPSMDCP37630DB5J6G3nVlZNn48gJ3Ik+gMWmbyq
oUMhkFRCcOw/OmrKiBH/nzp/DDes0JE7nyh3hBCa/0O0Ox9rKBfY7Ohpc5X/+7IDDrrRhE7M5hB/
2O+UHpVaACDEqw1/ehEab33lo3lXXV/ldUEJnI2HCM9GtMjjuPQrps2XJTtZ8z3H+0K2V8klhTF0
nXeyiJTUYhoFnCPmXqHsYskC2LXE0prpcHtOIXmupUekE1+KfWMTow0gicQL5qPAg0BjnUB/4H59
xKTbn7O+6I6ZF39oYWN40EmsgrwKkAPNMvpzUA9sQKj/PLT5Jo6o9iCS87NDB76ZTUBEe/VJj2SL
T6w8QXKD99iUNX751F7o9xDaedhsqNftVyn5pq+jBtQdFLnIJKcgLY06pJupWScy/V9fxRbDq46o
jleEVC+j+2fZZHnKalg9tDhvW0V9b+8llmSnw5H3y6ueSt0hybGT4ZIXiMsOc4QDSPs0lxrqI5zd
pO/N/tyYv/egpGPeLF17NhrGvJ5qOuikd+IZaqtCoCBXeF0QlcKcMmDaMIrs6QBJbxC8pBBusHVi
Y+qUXmEqj/AdtI2t9Vuj0viMqrd1WWM2TG1fIjqX7ndJkHEaQ48bVzk9dUe1+gMRTyf8ZRGlRNLM
YDQjUJwDJy+W/DrDfYglNtmg9NU+4jFJuRbuO8BAXUhrQR9742mMy41+Oux7xAxCgv8xe9EmzuQZ
vMCZdhPkVecdIB7PSyWPjnZQHIoMgod6HHDLHzDXWpwtsNZ6PUdsPf3iPlGSfaS8yxkdN7vybDaj
w9WdxIX7xtg6CbuS7x9iSCge0Bg4Je2l2gEDMiFD7TsTlE/+0lhIMSMIo+Ql9akUDJE8IB/lpfD5
1xkMCAWNwHjw8RmgfUVAQ3ULp3H2k4YPaVKd09Wm1fg2jV55BetaWVLu21cqsPfO1c8VomL2YaZ7
BbKAzWk36ICPJPtyg0W9Z637+KIztCjZhJDIsvkOywjLrWpi2ouZaAZY+ausrmusFvbFrkLynk0n
ysrP7jfrWqmsKjtconXQLdGzblDp5L+yJCj+pN4U/7Ml7bxIL8ZwQBU04CNo6BIrTVtGq/4oAs7n
64TXTWcrRfqo/ZRws6PeR/I8PVRDDfwXCujXi7ZtKCEQiLcjXi8Y18BYhq/KWgS74j802YW6uvWv
ULjPP6b9J+n2LsC6jpxkbZnRXmrWTdX9d7X1kde64KdvKjbHkx7Rdioom+7Wx6UJpPzxGrc50NvE
iQ3xtLWO463OX+Cy6mjdz67Ti9onAxmLYr8Vesp0ykBEm23nQP67O57GGdK75qkwiLQthVANT6E6
j/ungGvGVf+qzK5U7uk+N63lsWxjf5zRRCoXqgBo764xWf2t20fYnEvJn2CnkqVbB7LBuW9Ymq6F
fKu04Db1Urhh3i1wZC/Ntu4KUsq6T6jF5c9KjUPAzMp1eqB0It6/gnY8KsEO4S9q/sewrxsMXvTV
P6m0OS0wJ33Mo4ozTLBuNlbXjJb+u5AcwNC6X8MRe/OCVhIBb526df5ez8iSDu1OXxXkqBnqURZf
TZNtGwJ1vdIvbVeZrde3GhHrd+jCnDAlVpK27W5st/ioew67mjMOpSKdxrMmqYsy43BWrwFjlTFd
KjLn0bYdFUTF7KRYYTujiGY3k1p0Qhpq3a8YZ4++gwN8QiKtE4GW3AyfLX2xjj4Ft9Mv/ULhuvx3
voqfkwfmmTPm3LI9qRR3/rrOPjbZtMs73IK9dd97ZFrhqrGCv6jpBzKEC2Dojrqe01W85CZvwsEA
sjI9hv2SlzNIcvvrSl/gpCCxr97BbNyLoupXl9BpMIfv/QoNa9CuF5XzXi+tW6/QWRIh/2Jv12Xm
YOyxy5c+hMgB8BQ+yRy511a/6zgbK4c+ATZM9oKjXfjRRaqdgeFsAyENEoQfqrKu6rlv9tzBCg98
cjVixHW0muQOh/KzIhECIl2P/sSi+YTwWEqgTNUBf1PWlphPqcjtJhIagWFDKiz3KhDCpJIOnZ5t
z5WADmtkhqdc9KU1irIdUkdbvG0pTtVuJHSh7d/ubXicbzU8OYkFNrTawGTBFbfQg08o2HEJ3bgT
gYOpPDxeKUT0YGKtTSeObhk0thE5Jv/wNsmQCDLRGr/T4G/cM9ZZocSqd6HHNkRAWOQhQhSXbQRt
NlVwnlx2hSExfQRMbSZ4OP+1iHa2s+9Jfy59+7zkDqISzda8LtwRkdiWop/Hm2k2vfVM+hn5HFu3
drwChcvfj5Te5UNDXeLAOIOWp8T5oT0YdrhGef4Hoacko3JP5z5xMr66wP4ci+SwuFF5h2mZxMwy
d6YRmIYtLVjghnqiuIj6UGD8yu/WpLznCheQflmFX7fryo8aqH/qXKSR3/YZwk52/uuh43jCEfgk
a9NA23RFGaPps84nR+cyxIJOOHPIAvf2wlKmK1WVJNu9olhghsjK0B5GxzHD6hSZViRGVpO+xK7w
bWdJCEdlKR1cjxdIxr238lSgCocVnXYo6kY0WbPy4sferthPUMfLLXsstIjNaXIXGEL3bN57YmHB
BqHn4sTG6BsoCg9a0ZbIORrBM+EAG/8elKXB2z5oOW7rW7qjL8oSFcEuVMGYlXUEdyWIEZdekFkc
zHPT1q+VbSy9UaWpGFwx0HQarU70yOFzzYvaAUZgxCLhJVmeKbDV41YlZoUtDSG0/i8nvBJvLB9+
0DmItCyJnciABWe76C230gmVoTjD4tyEzcrDOy2Vg4dkFVrBjoprEL4FFnOtJRD5AhgndOd93xxZ
NxpCpUaYIIFYsyNtGxYg/7VgDIuCPjuchKI8p6Hr1pkKM65WuU0XWh3YKO6ESoEkWH5zdDiqiIqf
ZZdyRQo1M88+Clux4aouB8fb6Y4OZn+S5+vTWbnj49/BNXZX1mj1mA4HTk8NI+FAz9WfIAiD8lye
SbJEbRDcdwO1/Z962abgzgNOB8C24M9Uiibv24794yZKSAS0tkqQ4BnnDc4Uqu8TICebH5j2qLeC
sGIqik5VEocbJWNPG1mH/tjzahzxYH1PmgIKUTOVfiHhVUtA74uECIr5zqXuo3ETQP9hhO/y/lCL
ek6T2kBLVbnfwRkas4marCXNZGbEknIi1tUcwY3HoyQ/i6hKYFudrG4tKX0xccpdzssFZuWWHtAc
lygXwihkg3Fwfto/r54nZoeTQ3YElFcmlTr3QgIfjDH4U29CCdDZZ3F8vLVjhsg2OWbe1Yd9FYt2
jTBR1ps8hdDPoERWQ0ZBX4xOOS63UyUdBnVCWmimZoQLXLiT3k5L8JQ0q5MuEa4FmuR28Rs8AZwy
8fzQ4n76L6BXvODY5w0Bs9D+qIDEIba6jj9L+c3t9X/WI3CDmpYRVfA6wjGzChkXfH+UegYVUZCH
uBRSw5+ekDyx8/bRfHZpCUcLimJmHQVIG/JlZKQuyuq7u75qbnSgeDuAB6aYF2qiIzexMaOs4cAz
7cmb7fkbgk3PnFaj3GP5UJK304S9Sbuw7A2lgMNb2q7Us0vXUBIyi3s/Ua49qa+3v8NoFay3IrrZ
vEisqXzQSMXmvxrntLM5U/98Jg4RB2EpZp5vzibL5Vgy1XgSVAfFkUOo2HdFpcN5ssDdaulizPXr
/TM9j/NcO8ixRdm7ysJX+TCsnHBnPxEa0GuKOOOd6fLY/L5cMNmD+1jpEZArbfUD7HK4FdFt7RWZ
oM70EqWxkr72SwaFnAlOThbpJJ2o3wGW/7V3XO6vP6SaFbf9OWS9/dCPFRSGnrtSzMmf+5Pu1XVg
q8jvkR1tLminws2xZ4pv69JiQeF0u89Ai0Et9QMS+NZAPWiaXkVWkVeH+DTBrEO73ici07CIJpgp
OBqLwZXGMsz0nur4PGhbRP8oxGE+NM8O8CbGG9IyoglKHlWusF7NFFZSVCCVemIBA2RTOqL9x6Ug
MRxFoQSz6KKC3OtzDUTbQr45kBjgZFNSHTi/EB/zM/gJ7BuIunMqzA3AiJObMBsmL2aKy14Uqdbq
BZ91a4ro/58vVck3f8Zfcm4241jNTZkgQD+x9qZi9HLk7qqB14xiv1Y/Pt/hsj/oYF1Z1mbiyaA8
GbwLsk8k6di+o9wJT8IssQhttAqeIvXenEguJ+na+QROxFbH0SgceumOyGqSH/cdHXdVNZ5wJU8N
J6MSlC+f6+M5a2zb3nSxQbcJow+hxHLWXfRJH56a4GOMQ849E9YBJle14Izzn+p/InKI0Q2nOaKj
bTjJcHZ58887fhsuyC0fLAkkvZBobxDCQ+CpmuZ7yNYLYQLnp38ZbBSgu8QPpRy5ORq+JadcyzyV
1O/PCbGdBW1GXYhjjZGuKScRvtrJ6AA4rQ39DZERJkxL3qbiOVoigvP4VLFi5rcpJSbKZEIDiEp/
NY5Ss/ywRNPqp5OsgT8e3kXItDcLnuDstNbmA+BPDKa68lEG8G0Wh0ATP0jZVU3DcBv4S4JyP1Ui
a6E0xL4ugnrMgorRfQ/59YnUzjdsno48945JwQcFmRQr8QImEnpJcQ5A7xPYXlij1mDfGhA0O0TR
ZgQiDw83Tn6T/mUEr/4Y4Q0rokMEVqpdNsV/EHY9Xg+6E6nCTm44VaDU4X5IGQ+mJR8lDywCkL70
2t0lW7sxZ2UKkwAIeL9tSsX58RrX/KF4KlAnhG5JE7faOBOYxXBbiQ5/G0HvfDtm8XED0QZ23b/n
HYhvVgcs4YwWtt0/zHap4b6INqEMEpL2b0SA0utX0SMZZfVnHBVKCqy1abenUeVLSb2ITMdHIJJE
BQ0NKtwtgPtgvAqvwITBF/lul6swV9p5o8gXsBOLwFbHWYUHsPkPwkO5Kkoi6mIDJiJDkSvym/UL
9CQC3e7toMWfQKpiDdWBJ/NIoDxmmXVGlCaMbJZxBJHUnp43vDJ8uz2SvGZyNagSY32dWMvYatsS
jOliemYGuaAhhaY51ruLQE730ODMuY2C6njRh2O4jG3K2wa4MIcs24d3NIdBOte0kQFfFWaAbNia
NrqCDmwCXDxMA7PwvgrGy9u2XlTwCq9SXldK0uVUe4P59C5+qoCCZTAbMjmMi28ixRgKnJR38ZxQ
5K6uUllk7m+EJi1pdsyrKvVdfW+BJSvy0Ze2BmkSZFRMG6NPWwNhgUFGxgQcFGp9d7c4Se4iJy+j
0+tQrMudyzQTquT6VRa/HOAwMzVY/iJpDIsRkTouxXfSGiU7/44kPvZVntPWh/Lc5jTRWEGm/qVg
r8p7mn0lk4PLdYRo5UPZFbHucRjZpUWkhC0WqFnub6IBAe6vDzsxYzKtvi8v0huINGzgpmzzHuWg
xopeLkLwg7HRWdYhrTcU9vzm06FzP3QG9jSc/lPwE4UrtF+u8LeFCPKlSnMN7qi7Oq4ADdPCcomG
IEtulhzSFIQMKdGau4Itnw0DlB60E2xbCMeP8cWLbiRRu7fxB44ogw0azLjAe/DLAPRjpwn/8V7n
5E/sO5Lsibrr4WZvWHgYJ70hwi1VRSQR0iSilL1vo51/WeThSHqSOMB+dJMP5k9TCtK4sVaZwTud
4eZIUYz2BOLdk5KkP62aj329mX16xG1VT7/ywJKiWocuIMMsD7gM3wwoFF+e7ikmKREBB1mlAmS+
PBLlYI1nnewHgZL4zgPwe21Q+cK+JB3ebHn0BV1hzR4yz3AD45Mmw1/5G7s7euwiD4rRe4gnv4eW
pE0wKxMArDH9q7dcZEFtURtwOGIlo8W+QQcf5ZaZGE2Mj+PfAZbKpzxI6j0E3ihoMdkXfpKXxh8f
ryPcvJbBkrqi/lS4P8GhnM4vkUbB8GzAhpFNWfhyk7Nd9L/dZCzSkWYFgKtF3oFrzEvomAj8OEKL
LXWMzbysNWthzWLe6TwTwAZhZ2YxQpJWOeneZAUxJAWR8niJcg/PuMa979lJOw6BD2iE/Kjm3t1P
SMT4yedw4jxLJ3T2GZ3xJ9i5L8vrsNRDXe7VXI8IOVvxVHGF0bR476w72lJlmq6KB1UgLlfSw611
ostMMa67O7Z/RF8wIonFforcSRwg/WS/TsVZr+sEMy8YjvVLCIxcLzALvTTsosUm8c3gaYh3sYW8
+uJLwEcIfNdIsIPj818by9hRh2HGDB5c3VaMSPKt564SPBMkmUYuQ9iN5+Ro0drbmzi3bqCQVz3d
0g8PSqZMuyVNdOptQ9QXKuMsTZtivrrNfHXli2+zDSbyvMMENBEinl9tk5kJ+2HNWNugCq0KqTvU
vLK5RTYNEhpSOlGZFhWfOs2rk4sINoV2hLSzpLORSL7jDcmNoRdthUL/Nvdy94iWF8NqhdlCPpAu
czy0HOeUvhYaqCXK2T8Kkci9s45RjmIudJOoPwj5gcTR8NS8EOwLkju3FSOTNN2fgXhzs4RHf9YH
x4vEJgocg+FcGi76weVPzzZN8rBCQzIA4/s/bAnajzLxXT1fd98PbakiohNXs9RghXOH0VKugBVa
V+eZrlli/ufWDTznhmvzkx9y1oyWWrA8gmqr9jVa23+GjJ9J0jEe7fxdlonjys1kzBpThxA6NYFC
vjfB0R4+27/3HHKCq75feOMfBNUwxb4GNVcVgoLdHZRng3Fbcj8W3AreytymXMSG/GOKj9eGwV4C
hndgDkA1s8Qkky6YmbjQKtJIiCTRVeASQYxx+r2/WAhE12V4aohHQWT7evU6aouViFHQu82YMXbA
A6sJRWpxJoytEYfpzEkX5r4q7IFP90pdusZY7NvimCgVn6hHX+klhIUKHkonl6Jbz/ClC10tuJOF
0RXxXPusQKNEVtis3BUnEKbWjdgqjjFOxuvGMLXhOTZKS8kqEqEpl1YY4AE7UjU3HB0W8odiQvi1
SjBWIAfJJr5uF1In9KPMUqUQ+/1Re4WuRsPSEUtzDy0Pua7v5csV8LTs8VWYmECF9fRNPWWA9Qlb
y6P+Zs451N64i2wBkrXif8mscPMADJFeXL/7UmYNs9vBC9vWP00Wcv20Vh8319oCq7UwafRyOdlH
sy98DpYPCEMBZbexBwTKjhYJtt+qsgb0Cn4U7mr4EqNObQL7bDDWf+vzQmLphIK8Cv1ID7vN91qO
KI38eBNljzFoBvjh8HuGKyc27uIVDBS0zvN79Q0hhfeMjecP4C5br5+VLqSbQXSwGC2whCOMnOdN
Jch362LEYbTgk1N7TDqnoDpSZi9yziaP5hisx0Li42AqxIK012zGtkK3ozXfjsQCxzXDj00Dgbpt
8WUfJp6+v8a52X1FlHUELJBxzjJR1UTfAv5K3MS1fY/hkr6opo1aG6i2Wq+/1quEXQtVpU4+p/ln
xrAXCl40AUrcBhrd4jfUe/PcgoDUFgorsy7kCbIbTy+RX0xXHU9o2va0QtVRqm6VXFo/r7tAb56s
FpqYwNCjGvSFK1Db7HyUmPCaGidSAXbXfogUTZGDGGfYO0u3GK5/VvZDnYLahUSNwH9xi6TgSkJG
pXo+uDTLpwIUOp77WWD9uzWHxfY95KoC/048WZanb/HYrqSjhWJgJexR5Rnc0+HkVzGhUDg29y79
k+H7SvNlTxbbsfBBc8Cq6Kq0XIVcr8AMR1thbsYkjEhr0FJMLO1nfB9nXW5MxerPghMZkZzk3SFt
s63UDQ30mIa7sMkGUxG8326ZVGmQTrT23mK0XTLiBdRUHq/p8pLBesREdfSbElGXJgxBMd2DH99D
n/oS3/WXE5amWeAiAlwO6BQ9puJp42gfgQZtrVzDoIro7P/ZalWA7fQg1l2E01MpQ4GCYRZXZ1DG
4VY+CeRrkFzYWp37fSjMCHym8OK9xrnO/bzpEkXiNW8iBya3sdplkCdiDrniXPzpW+AyxvJmVFET
PQClpmAdAuj/YpnpyooUzepK4tqN+6abvRl0A20wK7ZaqwBmM7Sqeoi/DRIDgZikr8Iv/tuD4fFS
xhGUPYdgxFF4xRGFtvbNX5F/Br6cdOo7iPgX92hqNmWlls8IjmRUywR5AafjaYs1a2HX+0YJHt/j
SyVBAt2UNM/Cru6PCEFJXbBBCT88WmUehZck7xnrjV2CaWJknCWxxxJ2Gu8/oeaJBXWzcxXRX468
RFOPtZP93vNgkcB9lO+dRy/KfQxAKDuVrRFqBkPD18RfrS1l2HZ8PHPI38+cAR5/JD8dx28ig3QK
bQTSJcxKc2ZOl8VjhIZdO8mwXBBiwfhRsMat1dImdBhmWdgmq0b2klTOd43eDfwAh8IPYJ45iF/g
An6iT25FJ3OjWbKs31l4rFbwvEQzaNoTANG8wkjkWlaYM2lQrRhD4mLdajHlvCp54/LPQGCjLiiH
/yUo7y/vDDdmSJfBClEI5aIXA74a6gLGhqBAPMACQJODD28moo/juItuHZ0l5dlWe5oZZmmacX2E
TMXcr0vFNFLuxOJKMFfW0S8JGViz9Du/UizkQ/R3JKrWhR07Uo/UY8Phkdyr3+Rnzc1XONOGChGa
hsaHDG9YMyrR/ttRd/jYuEusp+CMh1DOPrkeIKX4FjAL1Un0aGBja8Mjc9u6UMUYz54k/ePU2fn4
VOrHTaH0l5oL9vBDIGand0TRC4/QlOCfcTnKCjDPLv5Pbu7eFFiZoMSAw6072BFOA5HFYMbys9wf
++TLnB3qmY3NERChtrCEXHTK84FQAW0ymvNSchM17xv0EYjnlnh1MFWFq08Mjv/LTQrNafx29tft
usItuY71dRZw2qsEEdAjdIMjgmS4ww0h9WEf9dRoD8XlqwKZNOQIV3jvJ18o0mzSxzUnfb1nDr3G
FX0Wjm2Y/kJ1Lm0slYQo1aHNho82WycJ3bsNEtHoscJpYPijzo9ibb4TzIGKwvQKp3jP4PlSg2XD
kHXcUmMXmtbxkTrEdRi77UA2o4PgN53CvYKhLDck+s50aWriz48mTIJy1MvlUpTFEjRLWQtdkzan
1YxYg9dtQwOo6ZCrPtwUqNRzCvtWfnyHsZMCYySfzMJWKEsdFSnPzgrvznIDlOWHRJ3YV2ir+GeT
ZtQYUHuBC4FiYxyYC2JB+w/WJS5NS0QITuZKJJPqujXEt25wjl/5yn4Zn+/NdNtVn56dGD/76vUr
Wia+fQsYpjterrF92xxuOLCgFmFWfwJKwqEZNz7oTKrTTObsP9zI6fSh3FPh7NLhjiWhOllxMZ2Y
XbSUCZS6JauGighdh9H7gnZNgA7a4U7xo6Yn2yGnlM5OShfYQ65P5k2v2NNeucGoLHY+xvfWUVnd
bEC2oWIgKlYCOui8a2Fa2r4RkHG3Ka7PGwznDgeB8yGz066VScXLvfiHNaB8M/gfT5QoqJgBQfoX
d1zwlOY/Q0SzGkeLJk4FWdWE19aIq83EQLEObDaKbwO/2aUlUO8uBkjEhye7LziFarZ/XYtbPU9c
Bd3hJAcDhzSBIHyQxLAC7dYIBF6LVV1nRljekzFNXP4SLluAtETcaRdjr6Ew46pXMNtgCsEY0dop
P/ALK1XunSScMwAc9yIJP4bi09I7hVwWCoqDmZGNkKmTZ7dsjtlq5J2FVp/l6L5IW5U3VnaHnNe0
lFo7+oz6SFNVJh2+/7dNzZ2myFft+Yc3nMbRE9CACao5mk8acfD//Pd+RSt53HpM01eMSiUy7pqG
UxNuM/aO5arihNiNR6nxfdnESltvqi+JHzQCPRdeFgEa6qyIsoVrV9OHaP8fMa/6sFKQ+XGanxzw
13h7NSPglhtOQQrDodBBPQzMNcjiOmreBUni6QOKGqOV+VSprben2PKixmbsyyrgvnE02qVualmQ
HVgmtVSHLHj+tLBNIXGvcNcsqPzqaEVCU/hsiDnlM8cBLQE8Ro0AU9NYzGTlKcsPSkIAzVLoQL5g
J1U0GSbgcKqB+v0kdhbqS1miWm96r5xzIJJXnjEC0t1eark/ver7FssfzpWrGlkDWQ6jJUu3J1l2
KTEeLi9Uvq7pgkKg2SHcGtfRIxeHpvo3xbWeY6cxOxsx09T2kitz0sNU+X7axuN9p02BLRzebUgm
Ei+Chg/louihJp7JcR613OJz0kLALHocMowMxphc4CeuxHPsc2NMHZq2/60PgQGbGZWv+awLN7ME
r9w1Mps/J6YttTmwQ+FS9D/RBzJq7cAQb6kKwHz2u2szCFc2pVFSv0Qn3lTFzwOq0TgXXjTiztpH
PRPHm/OjvWEA/1Yqyl3ImxaL2Rc71owmRqLsvkJegBZus6DG16SNkrnFTspiT/rYBXo0USI4GuzJ
lrow0KID2OPao55hfpTDA/zChcMI8FzHEjj0wIP4Y0Slqhq1JXypc4pmHvPMbz1eg7dpzvRuaVwX
UaNUf5zvzdRCoq07kcgal4m/KxG35sEXhs4LyOT6blhcfs4ZA3uMqMZ5qMgovZk/r01CozstEk1h
Lu55n38fK4ZNa7d82xfgN+KkkuX2eJXO5qHc1x+N3Daogy8iWwRew8o1ganAflABJksh3ZzjvEgn
GMMX5pqLqyP6EMg9Uufp8t74met6h/fYZy3SmZJEosAMjBVi5FkAt8/jYoKSF0nlSGAGHy6GRAYS
iJ8aylnelT7qFep1no5cLQP3JWDPOvZFwpaDVoJuezq1LFgLQUqtYQttJg3Ese9I7jistHttpiON
+SS6/PGxVsrACvgB0FLfvTp6MtYRiFHXIRO9JolyFJwsqQheAD5Yg8Dxn8olQJQGAMklBteyYQVI
yLCZsa/SyE1Wu85qc6La234Ra/Dtrg0FejSLdwh++O6o1GtUFpP0cIattK06AQ9HB86AXarb1oHx
iob6kEktTC8k7db+6/ZI9jSTZNu/dXmBPMaYtoRGbmJ48wtaGJeJNpMFY0d2A5h9syDQYUMjGYbG
ybGsvK4KSkKGkaW9FdbuStNLga/qE3JVqEeX943P3h6+HWqEibWtKiC3iaRkTyv3x9BxG8WSz0+z
sHfmcTr4IopRqfS7mscTy6rL0e4jHN0RhCjOYAjm0eO1sye5zqSw473aaZV2y7Rl9Xip38D83xTf
lovP72xN+vY7bvfJVjS3o1V1ICl/SLNUF01a2hhCrZysmsqQ9p3Mn9+AP8WykstJULyQcjpCnQF9
JMUaAW6K3hnu90KxCbihrikwYl5Py15GddUpRpGw+tsS2K21xr60uy6w4yOXd4PVLABTXHDAxyLz
bzTQl259MMPaCBX8o4FTPXplJI6bvQ3XkAyd5mF62/0yFkg0VH439uUNovea61QZz3CNRRkdFDr+
81FvU0XNPvVBwBYJKxXxGCfCgkiq30lanPxYp3GhsF8noTirwc9x16Snxy1Xr+GDiqSwt8aEfT9a
W6+ozoE92GLH2SKmCc6i0k3cu8765JnyPyLBifkEJl0zMHFeIWMr6bAIQSOnLvqD195eQ1iGENrQ
vxrCPQwxcY/A9tcObjmgkO95Ae9jIIZSG1ovbMp6d0h0Av042zzdmvpH4DPRuqM/KUsJdQecL8PB
Vi9H+CSneHP5ay16fqWf1qez73uQK8miQF8mzzfVp6pmGyaC6x4AKMGRrvxUC7V0JstegtaXR47/
SWCOPTRLhF2/RjE2Ka5/UPrJ+3/c99f40A17FD+o51dDS3CyLAofmdcPVVRjHqiyCvKp+9MfNRK8
maL78u0MP84Sdk4YhzRXbNOtAfggyT2aH/SmiSmKH5gJt+wkXWyOr2wV3V3LhHp7Os8zqBroiA/i
5HvwiEOnAuam9l+WiYWQ4Au+STcgAKaWLL5BcgBgtd2042WRanAd64k6QbgBYl6erwqE/DCHjy4V
xVheSJUm6bzWiMLIii+OOZiKCwx/gW9gypKDLX+WKhJrQOS0yRB7To9cXJYfaJYvqK3W+f+lQtwq
CEIGNWo12gtFXe98cj8GsLTLnOLdmsM/frmQeZ6bILZs+Co5dM1eZPnTlOMbJ7Y+U3qzBVS4beXU
TIkQ8RVWjBae97JrEOuFI5l77otWEmDskspKzdq4kqeLWBmcDc9KjZIvgtD8JSdix9C/p+FSYLuN
D1SzgUFp3/k3/Q1iOVr/oxAVBBg0BI8ujm0cix2GUDrID1AAT1y1JzRX1zKbj01VS/XVBMJBnTEB
o3egFolg039LZ46NMwdht3vY7PL7x6O1uQyoFWdr0lSZWT+dGsqKWCxU+rXgUak/Pv2nAdWP6m9n
d75c2RgGgqrfRT/+8FIAodqDKvN/sQq279pP6A3GfRWTUA3uovt+kFdZA3cF8+y8p84XYSdZcm1L
+kXbNElcuHKJRjUzGinZAYym9rvNV+eAx/rx0hZyPfFQud7wyHd5+/LdetoNHM4iZ+7TD2ZODaTr
amj4P513olnlNC0VIs36W13dPXA7PmvqdJPeOUCewSgiXn3nywQQclU42klr2phKSFYcXcbDZBIs
CDm9FA2HnrShXQTmCs8XaJ9fjueso7bXv0WW/11ho6rdeW3sk77JiZpRN2eSSoKvnTF99yN31J3N
+4LAI4taKe3bfmyu5o/eSM1MFHLzERuyzNU2k6ckFXezTGSIw6FEjQgormYD0jdQkxV5WxmGL2jN
rBF65DyIUK51xChHFZ3Gki7E1vfG3gag0xSS2aFjVYQJHKt9dAKDKxeqhQqZdX8s0glncAA0cXMk
W4I3mN1RG9Dgl/Rfdq//3H1unmVxnaXlWMZUpYA9UOt1t5FTRpsCLDE1xk2jhOfeXh0jRsH1V9Xr
oX/0nOPnrNYmnr+43aGxerlFsnXfTLb12bulG9a+YYkKRjbBIJKVJPJ0/bFdFhz4e46CMhrdhWSv
bm8hNfn1f1escLVMqFxa7x1XGoPxnOd/GQHuIsb5q7JVNoPdSJ7IvyneoeEze5+eCKCGR1RU1Pcy
prOVhNkLwEDns739F7EHqWnVe3kYHAbfV+V1Rojf2+wZMZWCriK3qpARvtywyszfPZOBdF5XFtzO
PqMF3rzd5jWG+TdgS+hoU5tttdFBTj7tlfBB9WHUtGKuonNk5Du7Z9uDw+bH3MPc2TwPTU9tuYow
IM+gv6VirgNy45Y6aCmdNly3p2Io3QqH7HK5mqCxRsICY49LZxgNgb6bdh+y3Cpcc3S6r4WnAFvB
bhnjIxc7MDyGkJgQQEXmdLfW+kxi9A4bEodaTHnwbPDfXLtb2AI+177gbNXmGv4x5K9jyTj00Yb5
X2PEFcSprczCekudkr1NIOfNHlM+/tvMxzVqd6TBYw/ET871nmywjcu+ZF9YLZGKlxhIXLc007Mu
tp8cRhAb/XMMl5P/IkRmr0UUa7Nlx85MNciuS6BpxkkPEwgn5jNylQlt9JTN6GWEmyQgjiyO56SI
HgOiJUuvN3xpGQo9sXjMlrpnie2386Gh1zqn7jq5T0PA/byWF7TdrEDlG7o+t98IIn3OP7P4LpMs
lOR5u7aUxQWn5F7cPK8HarSmF0FpWRxyGQzPHbjAtQvWlc/Dtbhl/GtYdcpKIDL4tbIEvfrxWGSd
38othgms8a7u2ctrlm26zmAdZOjgchBOH3POveRaw5ixTIQUKmjDDhvpDG9Dlo8YA2i0clCMKIbC
4Y6Gq6KYgVSOaWir25jgSkkvI058c+ZBErXPPg50gEYwGS032wRaGN3OnEga4CLzPEGBPU1bjFOb
xodj9+Lpp8HMkiPnjjSqSXXm0lZNI68z9Nwn3U7PMETgIa9fEth6JWXDdu5KUVSNb1OCCcar9PhT
YUwdhkx6Et1s5W3Kk7d+z2/FrTSZc3sWK7eQu+MQRtgCV7+F5M531dXQvP4C2Ln0PBivIvCAjCSV
D904wbj+W3H4LAn0ahZEkS01ORwoQAQuH5Vs9/ELaHwNcVx/+0vIZT2oUkMH/0T8e8jDQoaNIPPh
4KkyyCN3HJowUfkcp6ST5XdmHv1yAawXh39LgSDEh22TVYUYKWCxnW1xNaV9g/Q3rJqq26YLQdHP
SuvAd2MRxHPNh7uUlUSolU/dRGcLxHDdvihcRjEfuWtvnp9ouDzF5QV+BwKFlZXIckZR+flDo28U
kicURVZfyBd/aBl/j0XBJW6lIuzy69mUauZ6e5D95raZMMSaPYIZgTCR8VcWvgduzQXcB3PRGw0M
95RhdkxxEq8ueDWlBxngkO+rwdyEB5k8Z06znrPOChaNugpgpBfSzEE440OFbU7U7Bcfh+BDdPg4
AoXw0s83cujWMieSvp2zdHHlVJ7JEQv2OFQJBNi+AYh+nUtr2k/QZLpR4gK3C4pj1MUCl3/P6ONE
KmH3xTPPwDrRzXw5QnAQ0VXBAGNNlREI8jWx/0NHdlN2s95Npdggzxw0lkdjVopu/QfBckK8bFAv
qXz2cCIcQ/hX6V5TzKsyoM5+y+MOfM9Mj/8Mne8rKvQ0fIPovIPRfpT4xRjhKDY/VeydjO0v69D7
Zxbet+3fwaRqdA1S3IiYkyOfhoQCaPngwQSGJmTI4fpadvEZI6kYj2dNtZemEn6cled83Ekfc/yv
fUWoSxiUaQxzJ69Q4OTUpgDAkxu/fxgozNZQ5B/7yEZadQdliZzU5ili78LhTGvPYNXcbkNyIBkd
grLqTuqWk1nJo8d2RMSzivoa3TNKaHIWR/RKr7eusOuHNESUr4oREIfrXk0p+ZKI247ITJ3Bs83N
rzguhuTTA7xUDGrXcc68QtkWRn9Cvl5Ihsbq+FXdvrkM+Lmi4tHIsmSWk4dmN4iGox/CdFXqY6O9
dr2OubdKRZuhKtemMuCkHCGiSfF81Zf6FXjDlo/7W0Mx+IbOnu1BuDUTXx71K+nq7pIvd43mahca
biOIX8NsNsRCQFaOa09TCrjndny90bdN2H0LcJbK0gvUdNxRazyfREazV7ZFMe2m3ZmQFYTq/2re
NEiTpdI56k9ROTO/rWQHj1ME32Lgc3qz6UtXKAASIoOp0CZ38m22tZ71hN1A7tcQJkNJ2E1B7QNt
UlZQfZoRi71RWk+EHA3hznUFBYB7hNNG9LaFkaJi/X59rMydie2l5E1hVk5cZwnN2zndlxS8T/Bd
TQuA8EK8lwvhicl37Acv7ZTfJdCZRJoXjMD/S5+aeEQ92kx5HbgNEUAdLUXJcxOzRpxzDSROoN6A
IDMeKMdtRWo5tIhYuv4yONE6s+TZdXPk+UpcLA/gq9aOvSvJmWrhAz4EsJdVwr0XnHo6vsoCP61q
sER98u+oqb/BEITvo0AxzWj8A6He92kWbwpXO2wHN//xAaBwfo7ci0/YSD9D8x1enXHHeTrZuPRp
/qVab+FMBQWIJwJh395LaAKJSndenZTOvvtnpJVH41SFCOjwJLWTFlwHPhwVXVQnxukVhYyUgGkd
XLIuXBkmErz3H9s0yP9/bUAQeP9i+lEtuA6kF4VgBLj5ysh5yRM9sPrG0UhWwiFGS4d96NT0ExF6
vj+L39a67ziIwQhqvbOmkcGxWsnlBIoJDnxZlDAWI/hlnAQMoCGZg6V7Hw6VkHPD+7kfhUPxJhUo
V831J/Zsy3fBItGF8Eb0v6mBHM0YgFG+Gd66DVwcAY8+W6Z/b+zzfsdZyWiOP1+ItaQUKvZhjjm3
ybIBNQNKMTTF1uS57p27tCK8mACFOoCalSnQa4LbMUaJa/AbuN7V6sh7BzlTcLB3MYmcYux7NS6Q
0YOL3xx7EWc+EJi7RcYU45N/M1PIy9UzZqYIPlfgo2lFIV/AvcCN2b9Oi4ADGWmKEhs+fwxxscnV
Ya4rbJIeItf8z8ITvSM8n/psCg2FMnzd8ektx/YjHYGAGRH6TKvo1yNN5f6j/T1HafVLSTNW3smi
tbcIsAJP00D+4vmz120OHGTXtVgiGHYQvjCiiglvUYF/LdLjYJfghweZC0Tvu8PX9JWK07ngz85+
Ukt3useRPM6U5I+BgipRmZkJ3XytB596EucdbF0AWaBTLBRSTRrLFqgN3nB0M2/RoatL5NTsVC7L
Ipx1EmhQPLKX3SdwTrFpsElJBEm5iUW8mnuuZ9UGLJ93FqpsOkb8I4BZVIqlR2twtuKRXwFTmpSW
LMUOxZZu50vgFwyzTh4vy7uJzmrKZC34ALVhvuMnRoQkwr9L/GxJFwJqbRC5rwji6w9jW+o3qKp/
emTt361J6vE+zEqS5qapJ93a4D5rveA+JWEVztt3VO50bFtrAfsIj8mBNDwU8VqFjZe3Gex1eB1M
i2iMLFRyJYs/o5hFC5PNW7MKtUpNOeSsF6crHvmxf0VpfvUkGmohDe2YWKibA0eAttjdAecjc2+h
xT5J0PCcZOOk6iUNe8oyKTcmFhZ1pDgouwI8AhAPHEKy58qd2Xpe+Ill2kUiRs1MKmIqdmMN7c55
ChvJ6WAbvAMUK5bxVt/MoL69G1WCPe9D/Wmm1Na0f5eq69Ez8FF0zjKVOsPyyHrg3GYLP/lfYMis
SFzxm8a+bMyqbc6SugHhvwzAdLETzDtLdLGV7QtzpTv7eve5+SXLNcXd7rwYXzAUN3lcNpgAOiPD
w0dpeaSjyadCuK3FzoGVU1qlTgdZEJdszUxryjirGkH8IZ0fJ44Dy1PADgipha1zYo+lZmg1Yj94
DMATdvw9jD39NspuncPrZAtEHYR9vUySozH+3NugkZJTqmc9B7UY0zcf5EzEvekMdXsmu1DXMUTF
bD/UkG66wR9TLvqGZ/OD852JTHxZ4SxY5Y+0dU9LsqdEOcwSHutBg2XqUmbfTy9eOghld3hP/9Xc
+Cv58Kxdloh14RNuLDdsM2dZsVzbmGHaOezwu0Oa/Zq9YodFN1LlKDT4viG8InnBhrZ8UZJNMxR7
F1OjQP9hJrHzU9R0HQTeP/Dx/mHrwrNXRFLhUns04/W9VRFilXSpv4BsmFE3GRdPmlofYlHyaynL
STUK5W+kIfmn1J5x/Ty3xUbqPW3K+XanFToTH/nq8UPuJEe3mfaRJ7fb+7LK7IQ+RorXOjyz9cSf
YBgyd1z5k3sRuevIFaW9fNqzv0xD0RpYjAbGm/09an+LaUVvAAALmQodu9/tnRzTtLUMDG57fXaq
VtPauQ+fHxRRP5y/5R3zSXsQdBvDj4Q+cnCvIi9VlUrGI/6xq+3fXQi3g5oaA4NUP5PQBpOshvzf
hD0GSMS2NZV8bBLt6/EZuq0juAWPEAwfrYJtutjIlmUqecariLeQHXQU78rAiDryFvYolWzZoPO9
3lM/V570MZWS6q+ql6ZXqndxS7yVpohiXIOZLhabo7pobhvAyh6uu1rGDMtGJiz4OJEGgh/YA9U5
k5ml5cMxmk11amc8OWbwUp58tz2POm883c/S8u1Cf7mKkXUuwK/Kmim8Z5lbmkR5PtkpBxA+sNN3
gBLt7ob8Hb5L3JwZJqmtl2EkpZqBjEG3usDdXdLugeybRkm58qjkrKZhvLekYt4Wt6Lg1ld8oBeb
i3lbGtOjTcm6IqHxKBdy3PhokeI1k9h9fegTMhZKFjB8CH9f3zLEZpQ4f3G6u88XeFnRdR3pHALg
TfFkXe/b3zvnKuxC9WeDxcQxOjSI1j+MKRJwuWbMNSek/lNuMnDg4QU5BSVl11ATyQmzubl0gAED
jCzrb+GoXEjwGHAy974lW1ZK9Y1T9RaaUd+gN4HOs7/q/Hgd+H+zP5/FeQM4UNuI4gU3EAny4o1A
GxdQ5H4gDpfhGloYFBQ9pQy/HsYYm7OAUjeBKwu+W8GTiM9lonG172ghRJKQ3YR/lEqSs5af733w
aweKNIOpT/yC0RsO24XqO84FtINsG490pUvcHDG1tS7h84NKQrNJFLNOtlAPcKwRST18UdF79i7I
R97JGVrray3KxIFEXhfybKJnokLK1sFVztr6bwv16eo9JiMQiTuQCSNUzthsc+nsMjm+6CwljlSI
hgaZ/diipTuoqo7reXRbx4GtA8K890Fe2fmsXkFx95d0XM2/B0ehuJYSH50L5Dq06qqgUzl4D45K
0ptCuv2VGy/J86jlPVPCObcSfQVjTpK4Q/KD3J5JlR3PKNk85ysY282QHqfLP/knaUUpVC2YKIjF
bn4vVKB3vCIjDSminp2XJtDQOLqJUVQqYQcVCwxP6ajIgIBctWiNHPYdwkontoyv4BdyT/DdJH2s
uAdnHn78v8Y9aVzH8wR5iB8dqn1wIUKha08Lc7C24ETDntwLyaR43vPgRurz5YGWWfFP7JKKQWhY
76qjBOvgXV03M0CSuEwF3+zr2PyN2c0U4UOtnioKxxJrB/crSTFPj8JnSCuwzbRIQQBD9Fyi/3fF
jlinfixn8Js3cJBvqNfu+pl4fxhp38xTr2kLd73I8+ime3iU222O7EJNVVmtYVC4O5vGI1TEhu4J
/2wcrhg8xNGJYoXiYzgTCQV8eoWVXYfMhFI5vBMVqf3Jxy4as07mkjRWc3gzT3r66BxUNTOZhSNi
2jJnxK5CicXUGrVHk2ldRI+i+B/gYTc/6ACTmShjFrzFkuDZbWONfWba1W4uBlEmb6TrpOk1bnvY
U30ug6luRbY5vuxeXD+qrkQGWO5GLSqv0v1JFrHGIyFwdNU/+HbDFV9W+Oqh2fSQVZDhPh+nsJ/N
cSe54SVhGw02lRAlsEDh6jpT/cQLFfzzF2vS/VtQja9eSEDwsxYreBpFtCz3S9/ijpxSavZfSBfL
YkFcvXAIexPvZIQe4bt9Zj6weybMpIqsgGrHJdKVeTETwlns9h5OMhU73XHt3FaefTmWClXCgNIC
NFJ17Xb9ow/gMgGC2aev/m+lIvNnZJIsIwI8/P3ror4oPDN0bOPstQ7Tkf+nXYr8h6xXd6hw4zgU
1BuOWrGWGmCyOkm7h49xUHzySiHM2wEwHC1acNIGi0Kj1twW8HASsaqh/8GAhH4s9qvdLy71/pTZ
UpKSE7HrDRgVei3BH5BPywLb6GiUHwCtYI9xkaWivU7sWAECguZPvsoK2U4DaiKLiDEn0VW+F1Wd
kY1DaG+ulMeoy6HPtBGNZ4uo30knRniEQ8O7ys6rgTxtE/NANl2lUuljb734BN+yORFb2ZTngd0s
40RCJU3p5wxYn1gvw08e15zRTIR3LgGROYsJITEcF2j2OnHqc+fCYVhbmqs01zaVRIyCzQ3dgf0N
hD7C71vzvvI5MrrduIhTsVhrPAkTiPAsIKGlWmE3IGPz5mePMzu3A98hLYbwDsPCRI8578EBUUo8
7z36URkfDiww6sncunR0ZVTCPMglqitrM9BwCLs3GS0mSH7eYOOAhkD8z1hbusObUutUvdGkfl0p
E3iToOSjTXk0jWfkzGRV+xuRN295Puem/UNAcT/kKptAxQZXgTKxUJUr+XAB+Xs76cSq4JjCIOM2
CPo8fuNnH9MzIsOYqGsbDRgo4wodqKg9/YWdDyvtdL2FA8bSqpmCyTRusdV1Ws8r3sqkKuS06U+X
z0bWhGn9aokhOek8ppw5OjYSU1sdFquGsvF0W6Js4rD4kozO2rr0mj6uOqRXtIO7rfmGVOcPVl0X
V/rj9rHl1skdUqYgZg7iHvow1K2MvXJA6OZ3M1Vy7E1ohkVlUiYlODxhtvpcnbkBuid8AtCnO6CM
4J4th2AptEySQ4K1FS/OR8Jx3E/vvv14GFqeQ/HyJI9hF89vdu+Pur/kT4VWq8plJjbeRHSObT48
XE5QTPW2QWZAfSssA7L5CAOJlbW3AzvXrvVcbXenzJbHU3KGYEExqHJgn6VZW+EEps3CpYr+V4EJ
RMcWR+DHgCgagcJK6SMRoSsC3wjVO+/OtVzKuHBWmDQUxND+INRGbLazNEgP/L4ab2YmTRmOQ82o
fy84V3wPWFgfKBmAhSGLslQEexRxglT+Jpgjdbujkqi3Z+BUsXgFfDyJbb3DXrl12TUp9uqX4BFz
RUwawWjt+bXfQytrKglIbm+N5OeVgD+dE3mfWSBSSEVaQaYDHpUuTEzeVdksQhN9XxQyZBqXnRO9
l/LHGsr/bmQa46tQM+S+QCk/uQucFzP/QbUZaxFPD7haDsNAIpIRZm+XVWQJEjXzO5RCWBdGfWqw
w1fbz0frYnF8dzqO+TbLnipNOwDCITHrQNoGouuTf1jk53tglYoMFAGZwfAV477gpynDckeYAVSn
lsZlqklanreQssslyHNjDewSjFXhGYKs8hR90Z3aZW9NvWmtG1+zTRtdnbO1eA9ozpLOvpkaRREl
ee/cv49fpn3ojbd+lFNcyn0HbByy3hfifOFxd8fZ20r1DWJ2S4FqIaCJiToDspoxJVcN2im6rhPD
BXqHVALXhZP1R5TjEGcAwqrbyXsqr5eln/0Uj6B4A5sIFPdtxpvho1/B9PUD2PX3Cu4NUt0XS83s
bH+b9Tef8J66eRhGxKnWBhgv+OY+M49ue63FxZnjUvo9zU5EU888zjolhA8NHo3euhEupZ/dEPAy
rbkKc6h8BPuPUHYWFITigHYfm5Y6NCp/vq9a1WoGST4ovQ5rUZ2qmVs5sNDfZTuHqigkSUzKlp28
0Na5illp4TAKLoh2T8cpwgHRf/Nhr5ZAaZtInRFPU6JEXMK3Ys8J6RfgTwowAM7pIS6sOXTFU+5g
P8jq48cVPIghQAJCF4Zbun0PAuo4Ba0R8vOxf9tDnWibCgg5BKvRCwI6DJ6nUNCerqAeCLWJ9C3p
T6/fdDAjxyPovJfmbIpSXN8ZsFRMMChyL4XDMHXuCwN86AB24JDaBD+hqNPTZ100y78nehJ1T0Cd
LjMXSpniIFxv6Zi/0NipG0MMCmba9QioQ8LzXtoVCRdBx0DJlxeTuw4WWEi9wKcLJBigF4qCG8Qk
OQ2gYmLbyBbPf3hibzCfZBeIcWeR9sXvU4fIhFyumiqeLReUNh4GZJahACZ4eV54comygOrLcpT1
Tae7QRwvh5pNpxYIavov3f93kErydBy477SmmHjE/0s+lJ/h6DZv/HuQrmMAt0Z3U77UhHxc0csc
OsEiyCh8udrG7/sI1YTXEiHd7KJx9JTLKfdLBE3EJiv61CccNcg4/o/S2SK7bO+3EBiV27by1Jim
V62XT4hDcj859hUFYxJ/JV1EWT/Y3Ac6FCcm1StKVieYOCSWIYNBKFTbUGj3F2AGFNqofDy+VxRx
z5RERegI51nIg7S7qp08x+Km74lI/BctNdP9xgT4AlMwwo/ymQenn+nHAHX5Fd5RwrpUY4b2V3mq
SYUv3pAjRnUrimsvpzip5jNJggJDdFfHYwilQtirFdi5lt2B+rfZrN3zVHqkHnskeRT/WYIKNHME
YOPWKHBi6Tw+IWrdYlo53IOSPB1QbE/8z1FxxdktQA0dJuqyhWn5BO6AZFBYJ0Qgzw59LwR8Bghv
XD8If99lGHnvX/cfvnH/5MtFZ76ZWUy4b2s04iyho0LLp+wNgGVnQuB30lrRoG1LY79p/+WZzawL
E/V7wIJGmfbV3kOvc+4vsdheVA5/gW71SeoHflZZrgvshg7SUzicC1gq274ur1hT6pJt6ZCbo7BE
QI2mapE0JzIoqJugVe0UzLr+aKJoAviwbtYPk+v8ZTQ4kOvNtzCjUfd5TPNJaxslbmLJseiW2cxx
IkehSmhn3wIGEqvce86tNy7MvASCwuCMfISuySy3HcDWmM+QXuO/bpPoFNqNKvQluRXqmpvTwT+m
FcKPygIEiH57dhUqxRBDaAEmTL237kyp+1pYP7y0VbbLnIywlaeq7aHVLSdDWli31TF5GTkr5wtS
rpln3ltHF7TVNtL7WUMR+eurodNyE4wQscjYHMHR/g6Fv1FFVXMYr+n+ikLNM7iyhHF2kCl1ikC7
qCp038/2lDtEbMy73MBCS7N28QYgJm9R8sipzuxppkSlvmzCcpfpQNJFYez04rdh+Q4B4LVmTSXz
0OkELqEj8qJaklJoI//AhF2myJFGTM+41mK/9boPZJQfcaoNksMk9QsZm7u7Mn4KbiDPab4AIKTV
14FwA7onzR1jyrAnzsHq56b6wFuLBJFcF8tUtEpxAfAnwxdjLW/eGZOeGtoN+4DmtkBh87broDRD
ZIBrxtidpk1UeM+52qyFM0ot+IBAgvq5r5Vn/u8MS0pFi6HE50/m3evX0JThD6Y5n5OB3PW71EnV
fSU+r7aoogefQC2yvR3vPxW6X+vRonlgHWWlZ/FyqGTg3Vx058e5DcHVaFo+Ivo4aC7qug5bBTAU
hwUDsios8DLgYnVHjL15Fta4sX5MUTJF0q9Bd6/b5r1shDaofu8A83MTQ5re4d+3dS92BX4xisoa
QEpysyHQOey1k5J1ViRq7fZT+aqm7cNzD/y58uxEH4Ff3UA4hlftKg52ul/Nlcl5oEu1S0huDHMD
070vKKrl09G5+yk4FYie/9Zqz2i8yPJtNbXmIPCoKVHQzTprq5Jkk5sIeKGpWs+HaRXPLSQG3VAf
nObkeJxJmQH+JXuARdmO+ZQWwHLss9HObZbT4DPGThoLcxGh/K/PfJY/fhWp6dgVcQ+K/SdiO8zh
kFqC2lBkyf1C3eKL2YZvCihCo1lT5BNH5Kw/AiskDoEF+u/RvT3pqBayKAoFpsJAC685jyxkSRz/
qq+iAEVmzteMlVX5hYwB4YWFTm4+/hCC158FMsZim0ema+mhqoJoqP/zaHdCC0lGqXNBG46BKVkV
34jHzG0QbgxgE8NY++GWTKzckzGK/H0bhX3mD8G7Iq6hTmKDOXwpF5nwt5WjlhcNFqV48i5G0/IB
wtE/QnuXGuud8IQHkJy/OPfpbxAq12JdcSbrss9lkLcE4H356JadwEETOx6PVwpFj6pOJw/BqaLf
Yvqc192Pk75Q7MA8ykU1j96C1StFESe5MV8Mc18tvhcTPKYT9u0OKfZoFS+Ja8QfnLS0OJixEXR6
Ys0vENtK4MnS33B/AYzaxPZ2pRmGYJlGgfjp7Yg9phqLaS7091YIZMWpNZRORfJwSY3OAoWrCGjk
FweHwAEN56v7g9EaAiic5BofO0yj1QMgCl2knmyYhV8hjDbfn71vYir+YTMLkAf7Fz4c3MUuQe4B
ZWWS8ZJfVecwF/AYsH7E2NgfZdiAx0q8hEDybhYo0C1zl0pVA6qY9bzOg4mGb/oV8XNTmFCBIDSM
iXWW+Ys+f5kXr7uojnpm3SnY1O0uzcdzLkngsr60dxGKSmbDnnrG+L2gTH95NdUdQpTFWLUquf2e
uSUrrJJ3LJpwTsiam02K93IxZHaixg6X6YmP/SGp42CvOBL/VrzSi1OpnjMrWJ9d9FVfRLa3aSso
T3gNM8bEvxj2VZ1hwDE0CsxUa+BI0JHD291OO8eApo/ZrRn46hDsPDsVycJCNbYLWg3ffPuNrnuA
0jEIX8g9cUW866mZhW7nk+Y8pd6K+UDGmYRnUokWns6nTdfayr9WJx88DmTBzGNeFf006HDo0oNv
sxFP/TI6oLha14dMa8Qy9xkETHqeV+4DPh1SE6RMtbBPOyFMtn+21wLZWlPFiHW7/wAR/LqsZq7O
dJd8FOcAXR2mvf/s4m6T8XDxRUMZqg8u5ynhjh/voITukKfyKif9LaThjoNPI1OR9t4CcrSTdnwN
juaG6XRf5C/ZF7OlDpli4VpvATaUkl0ZvlAuGLndwpyLXFUZkf6rXfqqN221oE7fQMBMLq8mXVvP
odrcFPALbkyOmzuKgrh5qybpvF7cHQC/jEgkawEip/3q8YZ3w8yrow/Z+e10B1pvQWqY8uY7KksX
cwTK427wRFP4wfxiYOCMxtWkNtiMVjGgD0dXQNZEHtJ3OZWNm6jcTF6k/3ni7FL7mJb4QJKHKyOa
wcitaa80+BGTU9WcZ8F7ra02yJQjKc5bzEZRGBO6DEJVuI0aGAKREMUSasiBTKRx5DOU6TOfMovl
lKGM97W/4QJLS9yw/GBoPZbb6Y4dUXZ/cfUqJiRnxpP2yb+y4C/DfZ4uB50yqvv1k3R5iix/pIeo
k/bf7wf2vAlaGd9alB1vZ15BE8GTANgiPoE9yeBQGKfpdNL4rCVsSYr/7NosyMCHAmS7lOU3PWs8
OdhCwOZtIWw3x8Ra3gSp4jcYUzulvoWfbkvxE7LMZVXNnGghB9zs+bu7EiXDw+hq/K5ocdbQP3sP
4k50AjcYTFTPQC9Ob3kpOxHlwGVGo0U9/Z6SY2aq39zzkav6odCvrKnU/5sGcng1M4XfXCtuOrK0
yrp2g08q1lFLcCvYv0EFVPvdUuDsoaG9ZDBXiLjfP2XlhhHFxKGDDZ7vOCVerCa9ubiAPnb7usoj
UDzmht3CPkPaSAzUr6hXqHd4S9g46S7e5taaX+E/RSJt2mXyvd3xvSir7s71e1vkEv8wDpkNsUoS
AfEIbU3FjcAWmWdcKCtrWkaXz0zrbf/mxpd8UrTlAjwSV94hmdqyrOefx3/tSQyjZWE6DNkULZdl
xSayKae4A+a1CjjCKwMaKOZD2s4jUGPrlNeNcx18K7kcol2iwiOH350NS7ov2FhE+fJZ/epQIRp5
v4vv8HaeXAYhIDrD8uplSrwTiWmXqqH06/lxgAfZZTVU3nPxtpAgqphuQl1TMa7VrcL2wf9iBbv7
T1YuvVzio9jvgw1ZqchdMqhceqsh/MQz7U78MGbUPdNZaVzJt3qB3rger3U5OTmYp90IFIUInTbq
9jl/OnnWxModQGrSbvRGl5hoX5BZEeHHiZ1s8QmDHqMWpykCIoaWEKevjlq4v9lWX48+jmOxHaA4
tq+H5VGFK/nRYftWeXOVu41KIkDLAbUsMOZM9kgeWWdZTPLqrFCioYhev36ygWxGM2xIAEl4Orjd
U7mDaJAfPD/A69/9eKJDD0Z5CeDDi2IbkZuGzwYNie8IMugG996Mrg5+ZBiaHbjHp9ZSdiuiMFM/
SUkgxxZ2Xu5cW09l7Fd2/CkJvIss3xRcfC/Pgjon2Mc4zvNeizvlvw65yNBC8tFTtMB9jDSWIIcf
B9jARGbY8vhvQnNilUx4Dri/h06u5i7VbIAJSYRqUFJQl+s4jI3sfYR+4s70qq4tNgXBHDOBaa8P
tAwvpdaFIe6cCrI5DqcqCgNQmSqoet2D0Hdq6XNDSj/1UYq34F+2wdIaqmO/Tr1vHdbOWy4ogSub
Uye+PFkUTRB588ns14zrGanhd7YMm1P6tf8OsILb79jtQLCAKBJVja4MhVpLL5RAEdR7TMGq03q7
WG+BgHMb4MIjpROd662qLdbxOT2SYpeewcbx4AVkeKzHtykHuwEnLtfLzXa0CwsppGQjMthSqcdL
usloO8JO0v0MbGn4Hay+dQZeLbcipGzrj2IPTEqN29/FEMrH5uW5vAiZVl0PMaLMKkxfnSPMAy/8
82Y0WB3aGGHsDziQTDE3vlyKIkd4Kt7uYCdw0rXUsJhKQ4kEl2MMsordSe7IlCVWhMFGPxlcVxzf
QIvMgLkzpxv9IiVLClBT0lCXuQ5XDStbe3ZddVmGDxy6uzlHFvym+zcbWSltmyMYXnS/Cw03oxPS
j4NI+enXioMlku5HHeThfYcP0IJ1OafsDClac8eSs++HrbwPIiVYjpTmfIY4Wei0uUlUihmUET3X
Io1g+79UQR2C3ol8tQEshwaLUo5ItBPxXC/cJS41uSmbIfzFHbenz3V0oOrKv8SwznIFRGtMN0SN
VQHsX1EJ0vmrKAUL7+RfuS7OXzxyAvIdXJokaGiv9fepZM8hDGE/yz+EMcDI3jF9Gpyvld4kL6Pw
A8/Vlj4kTDCFtULPgCS5ja4Ist71Nq5oAkTcWwPZnG2KmRlPG71+GXUvfeUHOBfAnyrL12vC2ho/
5b18ExbMHkdSUs8AqIf6q5e5yKTpOm1LmOaKcy3uWCyaxcZkkQoM+hOTOWF9grBlPTT5DusBdvEm
eru0hFag/TT/uY5au/rR5voGjcVnnJ+8zNEsnBRfT8R+nbKwmmr2YYMniVuNRQ5tqMeKse18AQ+D
TatoCOKx6XHzma7E8pYk3EAyGZ7OHzXZUjpC4LZQxBZhd04zbNQHBmFhY+vuyX7O99J/Uv9ZH6JZ
YnNo8y3lONMJbboS/H0LIQ70OQZrHGuhhtp21NPM6qMYKXM7pqEiyUoQjBiOMNulZinHsMMptQv2
Yhrn+UG+gbPbkzoxjPJxAihYajqC/Kf+zdzxtKjx0mIVe/W9ZwaoQfrgr6YgFUPKXaFL7EBDrqtw
2aqRwH+GKvRWm6dLPOEss7jOGeYSRU9Lv5y2n6OJsIOk5YfGyTi8VuTggmIbhC7vggR30HuhUeq/
AuhsxFHwMAuGJ9Y3fk/tK2p9tlqVH7BtzBvcucGLLfhdjt40jyB4WjsW0CToztmHgOBkJjnwEyZz
wf1pW4J3Pe/ZUQppLMz+8b/w9qdH0xlA0ct8XTjRI46C98bSV3QIUtOIw36NEfCBIdykUu22Gggj
dpQ7RXxY6fVE4vekWI9mku60q8cqiNPZxCREJNkSq+eoolDDtnvlbNxokTbdNLL9o51/iNcvN4ZW
RMEUfrytLtf7y8i/91bBeLVVdTk4uA5b7INIvIQHq6Btug38+kyt21TzRboihYfq+G/4XRj67Cfk
3LtGFHbz8oOlLzP8BhaV2QbdwmkWALNycXW6WTTrmJrCDFRRx/fZsilScDc0h8JKA6KPCotp0CB2
DPh+900A9gFuDfJ54iSg2nmNqvktD9FA5pzHGy8yX9+SuCdQYkbFqwQqsBDqh3lWDZ0+lKmnRup6
S4yM0BK622zc2SzaguBt2LSpP17Rh/E9gZfX2jZBcPkZrYzgOJIBCPh4s6cFcZfpSFDeJtGBI2oE
uDBZez1TeV2rQZRALOgg389nT/ZIb+AM0T5gOtL4QgSxVOzfPMP3AB/ENSwMbQXa7hC8z6bT94ch
mAzBvoO7ylI8DUjBDwLqKqktMWSKOrQwEaxQUCbr17g+b5hsM5K9kVjenVGwJ9w12qQ2TjBx1VGF
Wr0ESeLhDdK3zsXNIMaGo/zt1rMx02cmXk1qGiePa4wQAPFIeqYCV/lAkNdPYdZ2wne8IDQFP50p
yYdWRmgG0OrlS4WcR86Gerb6GZ1rfdcMj7GeTOw9rzEZdfQpbN5P7NAkMXebZyvoNIson7lrVCyW
zovKFWbO0Wx4+BdaFHsJgzm8UTmXYwXQSI8LiKV2y+sf64UDv1FDBstlXqw1s0XmjkX1K9IZ4pcx
6OPBFsaz9JR85UA4KmcD3iAE4czKLn8GIr8kjBnrGtErxL4Xpx5zUa9wdRGvGpCVw5TRUfpR9rk6
KjqYoXJrowQcoBB4c6XlJRCYMHo2vLwjMX2Vsh0me6Vm7Z4HJ2cSv5y9ody4HCx/vMrcHxhuPXHV
gPmfkxW9C+StAno1XR0kqAH7snwLWmW4CLtg2uyIRBFk0SAsHhzck6PQx0kfYCyady9+xsKnc42N
gHYXwpMiw+nFnhp2BWJ7Ic8dpRTHG+Dem1SAAMydFiBJyLftmK7vNcSTH68NIx990Av1Dr+u4+ru
5HGsP3TvTNSO2AwSs5p4KVfFczDXcSCbzny76pS2jGhOW+T+0kDNebDt6EoCqqeeK52J9UidqZud
GcZXc1jumsPCd8yrHhcKNgZWXcWaBwxHbCGTMYipd/EUiIh0i9OrcZSvRf4PbvxJtsnH8efEptzP
EnEm5SWCfk7LfkeLcuopcnWvYQTBsCeWvSnJdeB7zMCfG1AA/rpwOtpQKIm2RxHXDwqcSAs1VXxC
ZoWwoN2/wZsIeUskucSHE/mwqXN4kawLpP39/X4oL/EWN6zPxVZrYH/Szb1ZhyHconM3OjGgDYtm
aJvPL0oGFQ+3NeVGbyJiowJXjXL5V39Iz8WXrM5iq+XqPscchtlR5xHEXw9IU6EDO4N0WVueR+o2
Uv8Bo4F7RPCsTmJBjEJH77N7z0ag6wUB9Nku95n8RJZEJcBlH73emsCCTBTwFbmy/XvAqX2kK+0J
beg31TeWQHuK9+y1kkYnKy6NS/cparvbhCng2VBzgt9/ivprt62k4uDIOotZa0JA01iuagtyvYzH
Tg6mrlvFmr47JKKj2kMrS9eH0WMycp/7V2H42QLGIx80EoAvqqS+ybZ9tbIsD4C5dYJrED89TZt+
EpY1sOJ62uSRckeqic49TVXLDPkUfg6/tXbflRE9cwQY+9LvnNN5g1+e8oLMMS7PSTwfnSXFb4bo
KqaO0lp8+di2UTMr8BgApcCk06JQL2u+Zrh8xnLHw0xnCU3+ZT6bWIQbZ62SL1becftvfT2JpXVf
QI5m3TGrLzQcEWRSPijEh5LEZirMQhi9nY+2wCST/VpkwJg7ZUOQVg0DD539ZSMeLrRuZCaFWcQ4
T1pg3s3KONO7ctHj+BD54ebjzVKa9LYYQFCXhvXG2VWnZZtgYvITPZIiEWXUUFa3l26npxD+YlUM
X+TUmJn1Zp3XPK1Eu36OSXYt4VyPVypMEFQCGm3DjdcbR8TQN2h6ffVTUJBT3Pp1LXkG5TtxW9XH
81BIdpGrkjmKIHGxqP/dLkLmxhhUEsaNOASWPRRKf0EZs5NbPIwXPtaqN/IoDWUa4LEwelAyvMB2
J5gPmZCf0IMBYqDR5eHK+0GlGimTztD62IdnEPZryihWXxXLXkUBL9Xg2QGdMHYmn4qLARQgGM/U
TEHeBf62OlusoqM6gnlwNFdWVTCiVJ0yCF8b4lnCWRHASWwUoLHhkHiYNZB3d7aeAu/ScaR1tC9Y
jdGj5qE5ai6mizVo2IEFZHdMhNAmvqjrbfBgvwMsxmqlk9sRPlQsBh+0KNu9IClZN/LED1b1d0Ad
t4edpCgiWoPN/td0++Occ0aIcgPYfXjaAx74+t+Co4sfwwKLrw8FCiEXjIlff2eVxe+sS3bFBxHG
TKy7j/sL3Bj75XrM8grG7RZW3V6vpnGg9rMs2tY43Kni5VUmJyPSlLOuZXwyaSkVMcezrb1dp+H8
cWAdXS9ebNkQeVYcIE7F6MVtfp5uKa3jW2Sm34aTRMnCrDi1+yivVFu0WJ6iRx5CaC9sy6k/VLjQ
NL3cXYQcuKA4JcNoTEqm7RYv50ixC9Zk1ZdFN+ErHpFr4cxx7gjXBsp8VBUQSW6p7PeONWoxJqBy
QDNg8wMqP5aAdO9oof/+HQYfOaYIkXhg4ie6sq7k8OZmnsQojMGc0j+10EtFvMk+YOHAp1AiOS0A
4V0F4qg9TwAr0oLsvB4xu4HgmTst1KDMJOBXjmW57MfXEVpivn3pW811K9V60hvNr9ffsObNEc9W
gdyZsJpaLUD1GmHvNO5xhfL8NQR0gM5YWz8pXXEj8Pani3w4jwKy7/+0l1Cfqcu0DRndchXCfPHe
6Mr8PDrzqMU/sjcTPDpaz+FhT1MjmUE4q2XruqRY+2tMJeAEe6sBbVceVvhhLnNCelGFDQzdPj8j
tCc4NZjJIaVksTTn3QK2KV0K+tkefN2mStZSMg+G2xeN36p9Lfs4o3bytRgEmqwU1pR57h9MBMZ+
tBJRYRgU9Ms3/b8AXC5sd1hqgETiasBNRNVvyjALCN7dRqNjetUjDfiGulepzmJQly2i4mQEgdzy
QmY3gWdu9Gjb6ysJe37bD0VTtCXpxs2s5Edx7EMLL/MTUCwpJfQQQ53YeTZpoleCMpwiRmtMo5xn
eDk8hLJX1+UjctgLubDzY4q+Caf79mWRU1auvQa5fXhTvHBp3wroFZIuTlWgkZrnjt9rIgYs//fT
46MtuzjI2xZdlL/r6+K1/VgnDEEHA4YXPi/6P69O7aVaQkKhdV7N45f8XgOsNYmSFA7Su74dmV+x
ZmRnt+LzaNTI73TUOfnjheQXMomxPUgZ3igej479aNEzl3lWvtvPfeeZT5ihEBiWS3/3U85oVlxG
54q+4Gvk42F0hI3fkIlDbULjMkhvkX9vFkfy0nZlKJbVut6CsNJrCR3dltd7r2Vp3UuD7ji+mxL3
MIRgWMCjv1u4jNf9C2oUP4ojLWKU2JGcvdhrhV3Lck5AbHby1+1We+jVkB75zFPnzDR/qHO62HYQ
oZP0PFyJ/fTHnQ8SMCysx9pWPA+xemo7uoAp9LRX5EhZuGhPxqWWTAJuLpzSS6skHiPSfrZYI0xL
IlGFjskkVetqVQmjRS2h85qT9PRY94JXAhCQu+ZAZ+cePbLp9xVaKHrZmfiDO9P94n9bm4ffmJbL
gay+PfGksm81A2YSE76a295FYs+zccH50+9U2H/NXBe+8e13y0ZcmweyWj6537ZTjaJpEpQX8CQg
gqwS18QEiMJ5GTCHZfBnPR369wAr6jIihWejO7RLmlwqpUgqcRyxdG1EbIKzuN47a4Chj7fvt3e9
iPTfTF7COysByu7bBNOo4b9U9HxxbCN0Cx6867BLEeoQoBAwlb4igzT+Jh0d+mBjxC1slC5pHI5U
xkIKsr2lklE1l2FJDLUhRGsOHPa//uH7xJUdjhMWvj11PdBxF0s4lZocaE00gC3T5c1w+xsj7lQV
cwgbEtphAvOq2daMPsNd53EvVF/psfWAc+89hoiX2dDYMjohrcXvhTlmjrdlNJK9W5afaMGjEFpL
TtIyOtiUpXMwPkiyipMC7Q2l+AUegECQkSCEPj3QsYf1lbl0SEW1rJrDOqtFWO4qToP2MDex8MQ5
ki0j/G7ZlBj4kcvUJSwzjqKDH+INHg3ZRQ6pKXlUtcKCyQ89KMjuKgpzwIYLQVGtTKqjZQLZxLyJ
WKA/jSuzgwjTQkREApUhHcYZz0pRYw6g2vqtUeS9XwUhUyczCt2n4t7/GJ+bAFmtfVawMC/BOMpN
jelI+0ABuHUm6fGz0Wo3HHYdHPfohApwgz1PbVfHqY8jmi6raMxkXRj9JXQlvhQkwG6xhEXSxbSv
RckoSZc0J//KGToHFlyDltJayZZPJoSfJy+mtdq4HtSEL7lU32z5V1vDwyhujfqhPrK6BEBKGHUc
jEcc9EwPvSvLX7SM6nO81egJceMFwhhXy/zmxuCfhxeeBKd8otFrQInorMmtAg076Xi7ViVy+9wB
TnIef0csXvSNI50BcEiVJYz9ZRsQQ7CczfVCoFGdhAllbfZXoLnyDNqE+K+wH2wvND1rOOL9LW2o
PvA6GE4+jppJ86It3YzFHgKh3DW+Bp+ObYKcFZxqbkY4IrZxemGnuTJBoOllLXEh79/9uN9oUb1E
uONewtqeUPeoKjoBiEM5pUxcr0ibgPEqPNGg9iBuXJd/KWlfD3hn3SxTqnNdrNllFoveXQ3TC/5M
k0mIjPNub4Y+Apnec/1MI9pfYdrmsKywiIMMthfiEZyYzLQWEx5A3Z46ve3Xj5DvJj/s8yjcbJZe
ESl/EjV6xWroBklpDfgqygUnwn/GNH0fJwPhCH41Nueq9SmDx8FbTLz+PbmpmOJlqc0jX1oFP02K
mv5C8uOlsR2imJUBurINoo74UC27xDbKGAhMEnhzunp2tUdQZappzGVROtnXyZj0UjMdDCltIh87
56fzxPhARhHCYCgwFu7WlV0X6wD6h3a7lPIHBWtPTTm8LAqWjGaR/EmpbTYGQxF/TjIrlrvMnM8/
Q2t/Ujo6ADkWNBQoTsraFY10Ny/x1yINCwE1NItZy9TQbvTdPHz9rzqwjFTO0PSbqIc0kdGuzalV
8onHGCd/QXeO52yZhvlWq+YR0stYJB4+FiVHvMFtkvX22AhoFtVreVwElBGC94jSiROrObW/wm91
1kI+hhR/gA3tWeto08yDDo/S6VI5uTPukAGkJiIrZz1ZKAkbnBW/Gn8yFGsX7dJ0s8IoegJ5qaQY
lbISvE3Qjyauf9yOrtMrOpF9xzE1d47yM0Aqk0IWSCnFjnxGEmy6hKIW1aVzaa1FDN5H27kaDKDM
xh8Hft2aW4RNIG1/ca76OEDNZRzK74Ef3K4Bx0Rh4FptQaD66sG2ot4dzfoWCiopBTKOULta484A
2KMMz8vXoUsKIBuHErquMYFml8+4op5DFeIa6BuCE6xS4le0tKgtctiIr/t/F3T6RXWhPPte3DbR
lSDh0CtLWSRFQymAzBgXcQHQPFD6m2gqGx8BqrPbtfKnFbnG6lmvIp1oNRfDjC2niur1Ak+H5L1L
knhnVNQviiuwS848E1sBd1saNSFHiyEwtmpJFyJulH1KvsRdS4cfI24UutWF4u2O4ogVeKJmcwPB
B05S+l1u6oBF80DO4ICpetapCWmOaLqXuKsIp7CvB3d7+qfnwVdYpFH075ykIcE81CQjUDAshYiS
opIC6mvEWdM/XtJjVPnuCgS/k/VtOYYm3Q3wD5IDHHKlhFAAQNfZP/urZjr5sBF3x5kUv5Gx7c6K
zrsU3oQy+UUWW+fHmEIgsklF3or1fYl0E07WNwuEQ3R1b9nMPt+nVkKVChGj9N2WRweFUgQPMbap
aHGWLhx3pg88c6qzTfcIbzkv8o4jVGbYivhjvtKqG9jOp0NpzypRgh0ZUAKM34f3A16wlKU71Kkj
93fff9oOi8LrLmiqvvp2dHozueTg/OPhA7xSIBTJejZDIuXaeoLMMhvcyQpyj6rz5bXstyNWRkFr
agTXN7oFVxZBWtLS807o8GouFPXoRAdGYD32qZieidHA7nqo4Zxci6Z2gRoMXvyBeVv3DH3x+Aig
yxWpPS/yQUv7Jvw4ZWamEsqETvrbwxF21iZEOAanqy5VNS8hoam9NS20PiEiU7t7t/JKlAzET2Eu
T7zNklNBozG9NMDss6A1neGF9x8j0IyzCros9PPopCrBlxpFbsqEXOaRPO6tM/3XmSc1BkafM90U
VJ/YmVYi061Sfsm0RQ7fOKUHmOrowl01TxsGuTha7iv42+mF9A60EGmZDicwq36bN+3YJ5w4slDY
lhX9RliTJX3vjbdIKWGvSUiH104kfRrP49ZFmVO1Cxnv5guZJxZy9dr+u3R9PapzdV+lJbIOEsv3
qfIS1eawIAcYvRbMH4MRoRk/p1fkuqjClkLHsWY7/rVz1HDtuL/pHvZ8L2OyJd7j32kjUZ8n3ian
937O/cJsa7GEs9k1Uz1fOsHqpUg38h3WblbfpBBwRhom+bCzCwXlx/laUBRVmyBDtkrJkNAn2SIu
18r9aKSYLnBAmHO69w2wWTk8jGB7uiVeoBsBUsSAI3Lo3kABxFkJUJDrO1tIJzHgv9DP1nJ0T9iD
Nk6DtPVqJckJq8amE7/X9/FcMw6OMI7B0543YZA1+E9LD9rmX3EslAgCMcpBshFy93wSB9sqX0au
2vUfRBFn+EBdNsnmYVIeTqh13XR1f7e+Qk1ofzClMkCVhDwDOXwFZMeuh90Xg8gGcLhz2BYzgVIC
+c4kWA/kpLgBxDcp9eWh3WyZA2M6Hnn7SVfFtyBN1p0i8WqQztsmrD4RylzUe1J9MTWyvmElyDgI
V0Ms2uyLyNTDwZ2n/mVfcN8VNf+G3c4sim1MECm3CoPrusL2zGuL40SX9SGOwmCzVdSnzmEytAhX
Iqku8384/GT//+JNY++uT5C0YPpnUkUuJFgAt0c1175fdAVpEPDP4cNxAAFfUyFytnzYZSe32Qpg
m/a3X9K65jF85gH34eAZLTfg5LmYl5d5IM/PV+IM/xnz0htIDGKyeIuFqzwmnQ9gaeRT1WYh/wbQ
RUCKdVWLQJNfQjiXVX1DuNrz6RgJ3tNWtql+kdTS39f1a/4rlrWgiuY5JZywPesVJlPBdyqpIOfL
52eu1rdBxBPuYvPls1TwctcvvEX/tWoVA0L//xWLWmhUe/71zLdrPc9+wPs8lhLqJv2RpoH8i6E2
jVTVoIk4RzR/k7BgYnUnqIVWhL4CfizAL9jHfVkoMth/zGC0Z/hGgnSmgOjt+luUlpC9/9wCRcrn
/YvAPGne6xv9VHo69940QWUH/Q0yb03uOTApOX+zS8dYveGPlikH7kcfSs2dsgRHG7p/1fwKi2p+
8ezdzhMQbD2P7tN9jeugDdE1kgjTGmjPb+7iBx5D8GTUu4KNJpk8RjVBt6O3qwf8k6rd0FbzF8KP
1UvagzhTVaEIuVxsB7emSxDVzwSV/bUXSJjoiY3uQIZm2QKl75TMZ83wbBS0HrTqkIKalEEReowA
iWRuHjbTXCq++Xt0zgtxQjsv1itTZ7TPFVV2iWGIUT0f5DOD/MoXaYv6Perm7rS8TaFggypBTapk
Nme/5b497YMKZ940kLiC+Z/ZZPIGcNCaKwtSkecFHGtdOXMUq7iWXrqNCuPUtNz/HNo9qB/7PKvm
EupQyZDoste+bxslTCoDUQMTKFk3cL0TzwjhVc55nRvYoYEgkkX7+yV/4jRIoq29n1XvdcMB/9yC
f4OyUT82Sj5Oxfn0+5NL4JXsqa3aKT9JSutfhQVw2yXqn5aL/kQxVLt6jahSY6T49x57pNPIPSO3
uNcZUPe6DhPN73YWhNVsvp53Sds3C3NsRTK1E8fR95YONIWS2GCD9uz7cDAMVDBtrT7JZr8CfXCJ
zYekKysbjMT6742dX9ojRVi9Y9BabxDl6O8Gy3bd5phyPjel3VemaGzE9u3ExUhaN2q7Tv54OcCK
boIb8Pbe6q2xphPFvBFlsCPKVf31IaCfv6YCTKMjh3YBDkGgoMhJkDA5rg3nCZGtCSegDZM8jwL7
Ii5jnZ26GQL4IpbujEAuHNR1Muk3Kr1Un7O2kS1Dqws1bQPlh/etTAM8v8R20IeOI8NLhaqFR7ig
SF0TcHihVtzFCD5feL2SRzGQ7fFjsYy+j0+ZKr0hpb6f2dKOt88+VZ3YwSCkZNF4yPsKUaLrHg/g
NhjVglfXXd0t1CArwp207WH+V8KzXr+PMXSfPfp9eaEqG98YapLXYSJvij7XrbdKw8tVx5MNqjoE
Vj1gF+CIsp1p5TNhlOe5iXhOKdF4dbpfI7UUay3yF3FVvq3NsQhBzeK0OdbP4bTP4K9+FsybSX6R
Dl3+qsLoW4PZIEZxzZzPmIH/oYb5JsP2d3+xxQauf8Z16BiAe8zX3e3J6oZm8c1ImtjCU7SY7EBv
eY94jryjwGnSOeMIjoQmf5yj1N0LYgqpCQPL8JL/p1SYtteSC7S10qj6bSHPFJCxtRc1Tx/rIgQs
+qRpsSzidXUudulPcPSVk+/Tty+yZusX6SCM/uHaKGGe2EErhB005Lruvo5IyZyTfI2tIti622mI
738/M7rVyHta0GWJ+Wrf1a1vmpCm1+H8ERj9vtWVSaMCQYObheZkiFhh6Xd+v3MgmL7r+YU5hUfa
ZHfNGDgboVHbukbzn3MnIRZIM3/MsmNtb45pKlTwRccCMffRYHUx6GUlBSKizt1PE4sYmrdsZdqO
7jwih/uB3L/XMFeq2EXl43JHMvGYUWYzf7AYdorMC4jox9/z9tIqNgITyZBJ+8Iup4AoYfV5QAXu
t/o8wHW0/49xsGoZYhQUywFGjepuhQJQALteY5x/eXwRXrXEjfLvZMIJ1do6PGV4kBN4DOFSeEGB
Iqki9zEWbuEQoAWBL9U/oZ2oBBWxJDCE47kjYFt+VOYwdeLXJL73FNwwayEZQSI6/lXFjfCFpvAo
GkHqUttmaaVAnx9ucTLQzF/FIEFl5WHBUC9/9L3y4JmnFDUgYhjhRIcDSv78Xyr+V4Vpz3NIHQM/
i05OU6kgVhfGCosRD3g82fytjLkKaVHcR6FzlMc5dqJb9eZJEfldErFs6b8yANcMLPobAl/mIzqH
gkWtzcMFTO7ixnBHkoNS7m21kLKdzm8yzySUCTfqXL6ZKoTLCofdHqNfpz3TsC434Sf/Xs7AwDpX
tRVtizXPCyVDKkB+2Lq/LMcEGkbG5bn7JpD0qqiES19ZWKrVIWLrJX4KpBgYMolN1XZimym8ZOxK
qcgyd0k80m6QH7ZG0FOIoNIElsGkFTiLRpsBONR4FbIFfEBSdxzTW2IRMjWCF9OLZnia7qtAhLZl
Beeu3ICuCH54tyHQnkxW9exVDO7LT7AkgceIXkginUi5h4gaChF8WisuOPludV9trGTC4ln3aSvq
jZjg2sCXdYP8qv1g4XfpssvYxsI9O8Zqj3seVN0f2PN3qZbKlJ7d6DAD9gKAYjGB/CHB7VUbsfIv
q5xypAOtnl6SzLZ3qOeY1ktvcnYUyUl1yyhRkJZoCSj1CCLkqVMjHv+LkaQCPmP5xSeGy9ch2vAs
+gKBlb8EYLM+sO79OrWv/P2+i0/OBbeHumjKs7ngSUJs9KVZuofBjI0q6nkwcdNnpKPrejqSQeGz
vmal/yZeQer3zPBUbMVIe9ULB+gb8VX7PpNof5UwbLNUbLwQs/s+M9KscwIMV27V8uckYQjgCeG1
MoJH34ejHliRd0KhP4kAyKlQWbqz1uAxB8icFsWodwTqF6urw8r8V+KQe3tMsD1fZfow0j/elJ3O
mHA76o8rrR9hogy+1XJklevgvVYYRBD7qYe/b1ivctFHs/8jOgB7D6GnsWRQMPkZ1IDPwFvG+slm
BlkVDInMVBGRS6E+0W+QCPmsgKHaWJC4oVLDlFJ12CZ0gn5W1q1yJZ+9N3zVtqaeHUjEageeVk4/
sZbk3FAR1tiHCf0L6oe6JwLegPiGh+KdXNX74SLOZXXPGxO8NnkgbkUOdA/QnmCDZS+Etid+Zadi
BlT4kQYxK5Eh8zjrt+2SutwTL6VY+FXVUutUrwy6oqTXKOfLR2xmVBD2Ub5lvY7GjpnwVO+4ts1g
YCd65UKuP/jruSY54iTUANObSMyxXTE8gUKogTYxr33Y7e7GWNSfo9OaJw3Av472TJkuDSI+YwWf
6x2QkL8kz2JgXACYFA0dcJZnqTLXJO4xsEvOo2xJnJU/Y1UdmRaaFhqIZ//xY8Sd82PAFq2bEBWg
SOaRY2vN6uk0j3zd74piFCSNzimyhY87WTyLKHOpZ50Z2D+3Xmf8weYXPWtKeZFsWMDGIr8irhwV
HPHnaaQW0iGxU4u2dyUHqab95EPtuSdioDtU4RKXpIjuD8cj9GyWabvAA0OCKWp9Pn4ZBnqAcIgT
PCAB13RnHaRzslr5KUJLgQ8HOm8ROE18NjN5kRJFCRBsbh97rwYbXwnk+G67h9B6j5b2YpFkW2nW
HP0fbJYeCg/QvoOl4AJ0WQ53+mt1B0ilGRfSiUv2ZHKPW4WN1rMmFif5XkNkGjLMllGB2Aiu3SaS
yxYu38rEXZiG4Iip6rmhIdzzOQuRFJBvi1VHmJOywfeoxajVrt/SgSge5CBvUvuOu9VrE/q3a4n1
eH+iZUZH3Wp8GeG/4gkEK+wTtD8ICHqYXhF6t1jWYjn4qUrbrdd33Yr16sPXXeQ9mCqeSC4n7+tD
vx+LUNxXKUxJfZYyTFIC/fvY7Wge5TSzPz9tzuKSmSR9owH0HBzy4UA+Gl/OjNGOtBvfwBLL29qf
pJVaF/jL2kCV3nLhodH3pcyTQzrWgJxrZjc1ACCsxGQEdUnqsocbo9cxOfsCCwcXxk/cG69ru5JQ
LUCV+l7yhEJO7/LcQDOanp+RohC2WRn0SIv0ofKCuwFsG+V8X5Bwqap1GncDlmZ+vFqGpw6LrrzM
N6aoK8fpno/pbxyJnUUEmu4ylTQ22+he1vySaD9/8TnLKzEOLe5CX0ak8Bf0fIqAG6zCgzIso6gV
Qt5Q7zOK5FxW132wEXqixnG03Xaa77X7RZ4aLLPgCvwJwIOMTbaW/snIsve40AMibtWfSrJZusDo
A6b0ibhQQf8SpIoRCE7IKii4j4fj9bj3jLTr+Znca6WvSnWMsVVSeDunqIIgqKOcl2NKff+6rDqo
OAPiBXhgPN41HrZeNGAytBStWdWT0NHUSWsVFSVHKKq6yUdYCla59wkVMu+5DewYTdkzZT0VHyHo
S4OgGv8TOcVrk6IVLYnoH5F143C0u44qEvuuhP6ANrXHbir3Co5H0OEuCAmoqf37dIU7DVHXr/hi
l2uDXv8nQVWeYOt6NXKsFYwi7N2AfJMZ+G0G0PdfmvDz5fnjM/+cWMCuIKY0zATlvW/x1og3sErv
NrNvSn9mUNdHRdbPh9JGd8Hh+9a6Gz1XscFT1u3yNflIrNy6oEXrHyi6nrJ9AHqA7o78xSCNoiZK
4hPk919/iKOdPb/pqyR8rJ/psf61HzQ8puLozq8j7TCdINFUELo3qOI6yFIZmORpXOv0VpJ3wtwQ
8JwGu7Te7PF0kuqFqTlYiGOn/X03Z/ggqVXagV+FMlcXyjUZ1Ce3hJwNUDEvt0iVNLgxpPXE/eUj
3gRW4O5QdzDyt7Cv+XSj9Nil6L99uX83Q40hVzh3xmM4c0WNrMRfvz54pmjKrJ//rENDOHpp3YMm
MxxQxcoNN5BtwRor6Q0CfqIuh/yoQ9TaLd9JXKFOYjEaz00EGqTTKBcDnT6aONwhQsHxQT0f4Nnl
fGpwFSsAkdeN3AdypmiaeJMTBKZ6Je9HS7MCec0FNfsAZmgU6gqV6ONvqYrkAXFN7Ik/O666JEOO
iTisCbMrbVB/I3s6I7WhViPjbygc0Sih1MNc/1ISXTQisC8iOAW8iR7ou/C2oFOc879oFXmCe2T4
n1gg9+JoJGmNcr4hVq4ZXtFDnonxQ69s0bizo37dHtXd7gI6MkU2YyEKoMyKrklF7l5R4MZHURwD
zlriqdQ+v+FeviZxS6BUGy9mNEC1oMMvdqOKKX0bUh4FAHusfdpzOpy6jZIEdhWHFXB9EW15YpEA
Qwggq99UtdNa4DeUF2ypnUQ68sVNZsQTtE/g6iYmwPo/dBAd79DqqIRb31DdwWG/M7IF5EadeclP
YUJRTqzhR3MPVlURReqMyobOEIgtoLznSuiuuaBzKk1/SZV+g48pAinlplGnBNbPCgRFQqjJfGEN
GII2r/ZxZZYAllQOQk6+0s8zIkZ0P/gZwrcEkE7k0zLxnyhoA9cED3Kp5wfghrXf2NVDo+lgC1Uu
SM8CbGJYsZrGwCdlsSKLDTFy3x4kg+/Qhzzv6QVY8H9iG5yYfy6YD7JnyvK4dV4qsDQs5XQJnh3M
lav8Vb7Uvf18IUmWcvXQDlWR3q8+d8BG4jm0gWiAY76V8iuea0Jw1HsYZAGhSrkRLcT4k74w/5tu
Te6EM2S14yDwYWoOdcmmVoMfegWVeMxvMyvuzMq0ywRmh4yScIpFUUrrX47YoipFV6FxgNyaDJH+
iCLwJzkjG400oHiY8e26Tdtz2t7SuFZylBTpAP0XjKAm9Vg13G6USUdyVe0fULFqhUNGFY0QT08L
oVmGtgAFSN1BbQmI03v/NcuhEa5gIgpKZcc2ASJlDZJuU0RoFofpGOTkcYMcSLmVAJAvtly15Kib
mhC0zPJL47/A3CdemOljGgXXBccSp8/UxiOBQ6TjIaqsZ3SV3+JO7th/Rq+WTQwE61oF2HD1DJPJ
8yl4mdso63wXwTMMCsv2kQE2DrozewBOdtXGFBaFQ3/fqbXLwHmw0s64u6jd/OsK3k6kzIoPL99E
xm++56jajmIrgEGHQLEAUKxWjA41+OD4foKFsixQutskH8KpJfmVk4wqysEJ8H1hVVVozwzeUOGv
ksRkqtBc1evhxLsuEf42B/sOzWtiOqfBM3XK2e0CxwnL56Q0QoyKAFxvZW7NRTQhi1KrzigJlJcX
PZ6iphWXVyYnwKC41+oGdkzawLbwFsn65oait+R91SrhTB++z+hJmX1LVtoZjnh3catEcufKMzcU
cjDkeFOhRPfo48IMjopNK7YBGRIE2LC1na4W2vQT+lEPcqEyrpmtf3XTitXY7EUhCEsHYfVDu+eG
jU6r1GdWxWcdxTk7dUoGm029PZ28o7EA/Jr9eRLYm3NmYcGSauC4CchLQJF7IvVmsdnE/FSUZ+Ns
Hh/a2/lP5ClD5X1nbNqqNU27RHfHCPuCkPEmd1NuyoZIcm3uiwrZwMfDwGS3IncnXipseqcPwFMP
NVxpOYqIQHEhiFFdIjSD3FeV+Eq37irrFzmnb+NCzzjGu8YIWBFZYpSWN6XXq7cq/5etjN5EIw+R
FiNQZm6BTxt3+zYniI5sqa7l9lAeQynd5VYucMNNwzVok9EvTOEoK5JqTiC6PNKonqISRlFWd0Ai
ujPsP5YhWapO8jVXcHTCS6i+uZqWC8IJHjg+A8uopcWwCpkto9bN6YzT4i17nrlp244fW0fLgVvh
R0ucO2DOR9RnDq4Up8AQc3W6DdjXzUCtiFO+31lZKxXWLu+9Eptchn8GbFCHke8z3TzC34+ppoBw
lNGn5xHB59dp0AyL15KlkaG7KbofgyrFm45r3fwttvhyOtADEsJ1JiyzqVIfPr+lxV6NZzBsMb13
nX+WKZKwR1EXGV0Kgx3HboUh6+s3+wGDCsrJMEcZgqk7gw16e+kH7yO+rmu66Z8SqwSFR9T+N9DC
dL+lZ5qYHDLpmxNj9DQc6q7KpI7KG4WKENIbwfBU6HBwUxMRK3wn0EypR+w3fGxto9UclTVYv8Sj
9Z76bjulSpWK5KeRjOM8QNPuYFiYCP02tD2rHlXq3xoSAdh/NhBKGML4jUGx+JoJyRnZrs99ISsc
Cvz5hAEmXRSlhWMM+d1ZeDMA2fkq7lGek2Fv3vppB0bfPqecijyQcl/Gm0R4bu6ZrWMg/fNOhJe3
VwkwK1EfOvvZsIvpJzp1E7KNCHNZAdZ9sF16ynsA3tPceufU/BRXJs+DxWvlEo3tvm7HYRQIx0AI
5R0PisdJ2z/06/MMSpHUdFLqdO3MNjL7p7XNff9TfWAC7Y1kyEi7lzh9CL/NCJjqVLk92bw7OxpT
7aUX0BigFz8SKc0z22lybq/3JYW3uAxYT1lO8oW+XTypT+9jNb+JkMyzosHAmKViGRfzLV3z/RCk
gF3ua9ZlecDw77PBeCZUBxZ2As00IyGwWmCDcEGlnx5FNMEVlylWqSXNWDYuBPW1e5pyzkQGOSm1
+/Q5ydioOYME7NsfO9wQMT40xdtYjjBbfM43G7z4CjSvbhy8gRocpFfrJMuCavgotkwWGSSROZAf
VbC34c6EK6IsmN72QGah0i5Fc5cPmniGSjUjx5VkeGbbiv3bgpM7cm57zYRySicNU8ixB0ZaVVIc
1QqG6uO01AhJG302qKIsXuisHKZGPayrlWFC6yus+gPF84NJ64kLihhm/bqV+hLfSXJHjgpHF1Sl
Fi6QvoNNaz8UfBX3Xh3DcNMhZCWI520Iuc4UY7GPNuUJfF+7+MJaJGijZDhHT4zcJTdV8EY35S7r
X4Q9B5xFbpVX5orUmfWebSzIYVScfrlf5tT5Ex7bQB+1ugG+HYRPRAzvwuaAXPClxCx6SBGPK6Uf
TwJWneJ0YoeQ0XXGsiQAPadq+OUzgp8lEuWBGEF4CFavqM7vU1zIcMzoqAbwZQCmoIe5Z75rwSBL
xUgNWny3xdEwuKUhDNkWreZUsOVF/+2YKMObd/oy1Vn1o7jeEMGGXIWApEbhXG2cYB8IOg7tdvNf
yu5CfTQsQANNz1JQuO/lxk6YZBvRzH3Gcw618belS5to1bekpUAxEVlgh9YOIfXi/JlVIEiint2O
qvRKlCHsLYqrxKCjV5g0Y8Ei7qjrMWYLrpM0fOv5BgytWc+SLYYpaLweD91ilhCvkxhylQF+BHyz
3Weeyf3x/6I+b22m089JvOPovTglyxfD5fsbsMvqnCLAqEDLODnsrUt5jwVEbcRQW0oW8Lh+GbaM
J9FOIafWCPGByPuNwNt7n3d1yzcANDY7WHFOQF58SQs5hVgm1jYRJ7C7/Bs0IsRBcKgtcXMCFOqs
coDQEjIgR8lroGKOGOIL2ufNjBj/6b35UY6hz9cKgpb56KcgZXTrkYEIbISMDTQy/A+RbKRTQbrJ
rK1rldkhCykHR8o2vM0bq2paOTLTwXCiZJXxqGr8LCFtrGDNj1rhuZ68jNNsUEkvjzPJZhTHwuiP
gaZM/4Ni6HIDte4OEoPEqL1zTeEmPlfXKmkCA0moxxUGEMLzUcAnr8UgGO0FPDQhJw7HUzUiBg7O
w7GaP+BjNhZPf2RdA0dLCg73abknO+5TFIHLjUL5O244CoL6AKd+o7Yq+TaI8GbRuuX79+sg1KZN
im29aB0QACmZ5PhHb6ILuddQq5XmWf80PZMRMOM/eOeMmgBnNzWIBSa4PI7vlrAD86vlI5SIktMg
qwybmV2Bpt6eSnESvTiZtFJysJP/1Ib/fzPxPhoBwazZ5SEcWakUwFi6Zt8XVsFSxmS6rbcwQS5U
HBQLWSa7QbySSAYgDXO11WyBpPQa1RZpb0PPZgpvzW5YjC7P1bDooeTL7kOlJgXcGLgFIBTyBqft
74ZK7yQQt42uENlzoGEBWkv5FoFVUGO+Fhc+4ZRZnrP04HZDzI/2XINcPvWdZrrn2x4Y7JJ/CTc1
dNJ51fTT+ouXAua4JWDoaKwbVeUVWlL05V7D9HrMJSZKLHX7zXhbUz2RiiwhbA1phEcHX32OvJIY
IASWgjhXA3G5gm3CjIDS8eIy4hT0S+F8UYejKpnFvrPRzFegcZucG5U+/ud3Grg2Ac2S5R7TG2KU
0FO+DfQEK1ZiD1X+eZ6IIbWniRLtzjtu5HWo3un8CkSJPhpDzqymeUCMe0yhnwJKOGPPHVoUhK0+
JcoKXrmT6R7921JkYJ6PF6pk5QxsAwywJyHo3quMBmcK3nlSILcqo7HhiYC9twQ+MDvmAbQg3FZW
YIbb3rSBZjuhchN72IdKu5Mpgbe1nGZ2hwWSsFkEk71rBs0UYIXh/3TlrMzf2ZggsjPiP1Z62jqS
VJnB2ZvvGvfxkIa7PYxFWZ7G7opDCulHq2QkiUkTcXRHYY9zqveW69mZ7iX/zvu1wRnhfDzdDrE/
nhA2P6dmApzdfn+riB9t7HUARKgUWhzlnVoiTCTk+ybQ2+oxBE/pQ72Tb/JfNd2nRX8pFQtZD57d
5DCDZjQ5Fm4rdV6M6hXNKIP2o2wEQ8wy5UZD1wxdkrPQOVWIUmWFJ9c/2uoWnGLjD18ZcyFU08sj
oP99sxcFgiIcGgtt2JAPW3vPh8KjlDNc+p8uL3ShBxloUIlH19i+KApqBZhvRPm6xnzUNEzIqZ0U
y/khkSm7ng4s8QxTW7bdGM9nMBJtF/+ctO4J6Y9HcSDtXc5LHaLGD+nGn6Gq3d5eJxGvlpc8T9UJ
H2m/9J1GWcFiklHgngsEb/rEptbtMr/ryTiCkPDEAF13a+AYgdQ/sSrr/d9rpqPthnUfj3eiy5i1
v0xlZqKlHnFqmz7dm83N7q/GcVrWCARTx23uC1w5/zIYna7VBDz3xeSBaYei4pcXp+Qy/U1IbshY
hY8pw+ra8X/pWOxqU582CMhWG5jstoI6qmEJGccDNrOJIctCOvFju6An6OKRnB8gzFE7Y/hVMvv/
BEuhycXFypYX8UuHcLJRxGDBGvpp6396RQ1QDQbnPmpI6Vs3KHi8wSWwuuMaYN48Xtqpy5S9sRlc
Rrg5OxGlyjC2lhWnuf/3R/lxcfL6NA3uHNp3jekEqb9ZNC9RWGc7AxQ+lbgmEpzvek4rb1dp3dbf
l+tHUA/SarLlUkBZVwVGXKAUFbhbKS40ba7n/r7VZZfnfG7R6YkWrqdgYfvDvpk8NZ7sFyJJ4uUm
kF0KjW1rZCWSxlVNNSIU7PWohqw2iid40GFkBKz17YA/gfCeaO1OqB2CroI2yB39or1YA13B1gxE
RqkYRlX0vy+95dX7vlYTUkR80Q3F6Cepo+RqgvcArd7J7gPKmUj8afOPUEX8JdkGDvPKbWhebNGW
9zGyV1yFxp7bv6C4kHw3slaLc4QUgem0O+Eb1eWLypgMlRUwhEfy7G/FqOlc/vwf6RUHIcSftRGJ
tMM0gD87ZGBFOvIkbn807e087AUhSXRqzYEQcPcjq+Jr3A2WJOqqbYmghwlq4SZ4cykzzGl1Zmrn
RhOAcTkgYdFF3q+nEdp86sIjcmfOxnwKkA2gLzHfFsOe+IYiuwighZywwTuBlyV2jRLafEU4zHUc
aZ+XZncEiII1RYJBGCjeCSYgkPOt38e3WMFW75MxqKqOfUiYiu9vbB3CSSLoZIfRWQ1tdMMNKGaD
TeEIoYH7ps6gZQ7ZdINO5o+ku1bVHn27UXsF7sL8FM2jGUsmZhF2ysJcnR03DYBw9KwJt84uK60u
2hmx8PVKktt8Rj5SyNkY7zNnNWy9c3nmhpI15aNbC3gLuL4doQ65RwIgP/H7QaCgk+53WSYQ5nQo
7kDs8AO7odwrFKSpUp+GySTmbQiFjewHJoc+i6C1RH8Tt4jbAHLh0WaPuWfMHIFAbDBtrrySCM2F
8xcVLS7YlzBA1RGhgEQJUrCts9AIFbOYYrn+O0EiyytIkLzLODbvulicD/jQxoPHcvNykoN3Qrdk
tyNtWxzeCcMs/qtaVymuSfwvPGWiXnWN4yXrvHC1qdfJn2grJigpE4sGxOksRUiDGbf2mwmmO2br
g9XOVLeN2t2pLE4VP80w8VVL75YxOCBjEVjK9JRmODISQQdSrMXBg/pwkwEzVkCLHHZHchSwyWo/
k+kMMx46I3DSX0+dWfr/gNM8LTLyAmAYCtR5pQYsIO52UVeZ56+TTJ19PeHfpNyHFV+GLoRMRyAO
eXHaRphL5Tx/R2pYHgc1SHBjYO1+Z1yaRaoTf8hvWDv1BzhPuFB/qlvZ3/SkjWeE3vAZv6+FVZYo
tPjgO9InJ4cJZys91JiTwWqYILzyPNYJY/mdJrKtz3nnBmjdq40gad3zgujrLPvlEsaLXNLqrUkm
EpI9biBBuwOz4CUUisnVXyF8ivwYmj83VsBk7vHIUdoEs6BaCEeiVV+SNgNLyZfZFEez1aKeAtcj
w6NSX5JBs5UrFaN/Frv7UfvB36EQf32Un1unZDFFsRSBV+wz6yrSEejMW5zb2GMHzaeeMSLtHA2O
6XDdn7pEwXJTOCvG7MvUxBubrNEiQL+vNdwWWw9cKKR01hKRiYCBttjVPmQ9GOkvuqTZOrL0jqAJ
APJMaprFeVmebhLoM5emPCnfKw4PSHzBie/x6cl7J1k1iIewm+ta8D0zonQ3Y1vmNVXLVcX/Dzy8
CctlsqJ8GoB/9zrfVm80SdyU6f5ksYztfXrpl4uHm8Hg/nmZLgrILdKbVy0j62qmffj51ulP5phy
qadxfJDtuNo1VqBg2cWs0+6iGOLn5N47UwzoCJXsnHUwUDCHISho9eKkPhcgz5KtNJAe279BhxxK
tVdJ8DuLM9PzFvFk4SyrNFBQ4sav8Hnn1GyTboXZdAdUUzAXlI9hxYXngFfYAk1RYDvdPGnYOLMy
4dxM+lkE/pkUW5smqlzDPn2L2702r70CPgg2T0rGS4G7AbA2YbOPCTMLrG+gGKkkzMl8L9TrVIwa
oE/8maoBBUnDQRNUKAqleorMkdTv/eaUJ/+9OcEFwgQ0o4w3AfxQZ075phPEy08no+eb/Tn713NR
xygsLlcKaQ2jFVDLxZ1L8Lcgg8geNbgOcmeoAKm/0txs0Vjhylj5HtxfSkt28KJHEXPbqgLaRguP
aPsNmu5a95waeg9bruFQO9he84zlk64V0EKTVN3SS0tA753cnFHUaF0nH2U0Uy0vGt2EPWI70O1Y
XeLdtKXU34MRyHTAOkVPfDKIaUDgOFaYvVrCYC2o7+irbcB6EIjtf6u2m5GcDiKGcQkTGhtuErg8
WObaAq87ewWkppXpqI4HkXR997fLPu+6e5v3d3J2GUp2ESD5msT5OsFJc5Yy7i+Y//QJMH9puu+H
r56QRwAt3sZ7jJOf/WS/qkCINcwElJADkCj71dwBRSRKgsqbDhKjfvLv08MzxB/8xIjLiaCOwprp
UJ2+4BMvl5tm8BSjSWfRGNINOVT3n7VmJNwgWyo7i8BEwrGVqndqEU9Bv8CrdXZHdglSpqSUT3gh
NBb9hirH7UeXBeIME3FY+Kr9LRhGdbMzRyOX25PIy0te6YQsMs5f/BzqDp30Z9pbZBBMwQq3RiSP
Y1VbAuVTYcO9e7XephPRs4x7pnO2pB0BCWnJIt/k6SbbQC5vIhqxAy8fX+rM1ANHfMbAnex1VNw8
OItp+Vj9X33r+4ZKDy6LjcFWYW+DrQePKAeaHYVqvXpTfu8R5iDTWVF1QHNURCnG1rfNKCAwkist
7JBHjFz6WYxuwqpNkBs8LbdUeIuy+cZ+8o0iUlGT0I1b4sMSF0Go4wNWTgBginLnz0lrROYPL6EK
CcuUQf+PvBWt1EaYgBxDTGv86dndh0Ewb98MuntGfBCsXcA7mL73FLR2Kn/efb4kPQjrarslztvn
PSHKssqPbPIAvVnUDuKspkm0EYghfFkgrqZDU55+uVXkQbTTUWwc/PfqZs+J1FmZzhSmsErO0ITP
67KO7Pw7d24187GkB7mghKbci0Zk+cZoG2evNRzAmE0myjzyi/oPz5ARBXN/ecSTsYg3j84bSuQa
uVYEy/iWL71CQFOzZyddVB5BeALmkhQGQY30/eR0Btw75DoKR1Xcq/y/Alljtg3SzGWu+qMIMQQi
pFsUacQPEyz2qBN/cXUJKtOvHs342cbJbNe1Gi2Fb7MGQYP6yab51C8M4pfxVHDzupAMt8Ufweha
7pGy1ZuWUfUTI7S56cf/0rIUQkqoeRJLS8gXd1BtJJ/ivgsURxeK3VISa1iUWpGFd2suPf1qYjnf
gA3aE3WNkcE8eIRxbUfc04hsS6v1lMrH4qp0MOjr+mM2y2+9vUX2/4B5sNJbYDDnIVA6le1Y8CVZ
RkWWUKjt/FGCVE0QEOJMyYtPATz9LY8fRLQoiaF7DVqoOitB9hiwQarA8yIi0MgBZueeYWFyjnAp
xX5bOrJ1lSSxXk+Z79ejT98Zw7IEiwxDG7+BtUbXJ+g5QB8AQuyslTW55/eXsFwkRrgd/h54IRQb
TxIHIxuj6sz1Ex/59nv0yZzB+4kaRH0iJTiovRQ5SsDVKcFNS5+XJAY4lFUBSfqalCqyT2znyE6r
MBnrAdDAruFWiFS7/vWMGoAGKNEXTOatP2IAKXGd6aljN9Rlc4sQ1p0LHn247ndSpCUKe1qIJ3nI
k25dOTveQaG1uwWpuD3dj8R0UaUEcNKhGkemydX8B8eQw6IRtKMgnv9+Re/gEH3yfrOjiiRA8CXc
6HNOEW88vCKg8ZxfUCYuKhZTrlc3G7pqP1ApfY4M6LhgSydL3XPWqx3x69TLEPNyRNJypwPRyWZ9
bTnfiQFocwaTY+lqPjA6ZimJzEIvz0i8xro1gNVtkN6mxoih0HBPuhNvouYZbdKL8ATCzsuaWZQw
OTIFNd1ErNC7/WnpZ+Pnj2g0FUDh3DwFTe2IvjtBKzhFRH/rzdjbykWODTMXKgqphOQoAeZS/668
51B6/tW0DvpJRemso/FKkPXdFExOfNZeQNETjCGMXdI90vrnXuDxSH7kaHkPy+Ors7JodKKn9g9R
ZpSqvog8YxWoFZaWHaiA/wTKU+rruoP3stVn++yDIu3syajEFKPqBWNFf7Ic3ckqW1qL84DUwdnz
1EY+bloKJGDjmM80ZSF60X2J9ae55VL8ZiafpNEVZL8w+Mf0Y3Wb1Q4JnrmMiAp8K9DaXvHf1KcM
DOmWlqgjL2iEUfOOhIhJDWKe1gcjlPUDzdwARDDImcBgkGrd0HRbNtcw+PFIUA6zWoBpCZBRCRCs
8WnKtyWq0Gc2Zs2g3Gb55e5rEtlPs6pI5uLRH7VskudWmjuPv+1JdCsob7bFSz6D4eW2aAI0rih0
WNEKW45EYmJWnQEdKXvo5osXECdh50lNWfxHVB4+2azejZnkBVIdtAbAHU4ji0JHqOBqxfrRcWcj
r+Peb80D1koe1vRwfiRLK38LfqpRHhzkaAcJvJSSVnNWsaAXWoUScj1bXqs5pkDIdZoDPE2vk459
7H93vP0fskHFtlBUzd1oYs2+8hR/H/3Cz2k72lwYomMiLv+tKAyvn9Vv7ZAhtq8PMhGMXCqssqs6
axY0DsKXTiURAmgZHszp76da0kxWRLYkG/6uMLBed6eB3qPEvqgw8DD/6IMQ8xKYzWGlpmPwMHrb
s4bN0bZoWaEd5urLvvgmimZ2LsyUPcZQdxC4yNgsIx2vZK4FxeqRdft9gSKJD0jT0laJ/avwC0O3
7ob3NdBFRc5693sMIphNuPsLg0SCHFDPK5M2+7sS5yBnygwlY9VJaT260NQjNt3txnvynsBEsp9/
u84xpWfKfzXfxQiaXv2cwb0/DokeFbeW6/IFyNn7W+OxxWUH4DZvSUS8Zd3XRFNII7992EPPZrn5
KJ8Pwha1KXB2a/MpCMOScexyxla8fZct07b6iVFqvpXME2xqw/mHmOJoblUdjvG1y+bORl+9bZJO
a1bz80u91qVgHrjA6bQeeqhMcgT+UNqPgReTPUHJH9PSM00VuVpONL7xLG2+hsI+zbc4548771dH
XO7zA+bRhqlBzB5BMKufNL2N9ti+PHJAQLldwgm3StqqDqZbrCMH73wz+mZ1e9WPeOw0EFu3vBqS
Qoj5VVaP+vdfqiJqx7nOdYhqJa8+NSon+v2s83oolHacIzy+GPw9RNDUu17DDdrMMDqWcPv63424
eHfHhVSKa6BmmZP0CdOA6nbVBG6AwhumyZRn4E6jPUFAlbr1+S69BVGZgfDXaH1Zp/J4KAPVwOtW
D1SnuJtUpmC3hk4IgXhoq/3Mh4Vy6wOo6WYuv06p0m55wQUfmSOcdM39dIHwJnWLwF3JeGxNNq4i
MXsI8oCP7/qxQNFzdU1USVXM6WmJEzg2WVp8i/c8PnM82sB67NlTlIFEAV2NW3P+HTsCWddpND1r
um5wO9KiYd0JbLBTf+nUZYfD6MrCSDQ1gv4Lrqaw/Z7/C5tC8FrMCUuAbwhI2N6Lij9qLzMIPkdy
67i8aGRX+aG2HKZ7dUpltNV22K4WOdlO8lRlM189xaP8D1vmMz+0Ttu/GOpgp3QFJMWLAKL8hchg
PAQsOKaE5gZcZONjy2+E++6ej/S5gLnG83uyiaDEeNX3d9sacfIAKxxAlR5o4mPHApc48YW9VptO
6zUVnxk7DKsjxAXPQ29Jl5rjbSHYJdoZ8V9E696XpipPKk9BE8uT2jTtTRZR6CW3u8cU8Fpe/L64
Vtm99320RYJ2z7m3vUs/O3yI1O2ignvYS7fbNMkNSjFOEK3z1I2F8I2tPo/2sW5DQRlh6zvGjvIr
AbFmkBU31lhw4UcqHbYP1sFxlfMvEqaTWDiEmGZ7aSY1MPojLQohWG+oeLHa9E9XVykBf4/XLtME
h7I31YsXcv2ibtg+WbiwTfAoFshcwdZUBiToJadMPrQDw2f4jogHhrH8ngIna6RrJ38TT1bmbkq5
emVGzolGBr7zBj+AtVdsx5vhZkPouyQkTWVUlwM/EUCNY5YOaoGflA8YTxoMEZr/7EqUyGAYABNB
v9Ac5RIJt6vbOigkgAewHvbjwcusNlXOWnNXj2OwvVolUSM34z093oFldcTxm9vJSy7AZ32PzL79
A6uavQjry+Y8Ur1Eb8u/jGpD92ZgWu/SZCMtHXUDD00N4XftsN8iq7bzKioC3jZiNaQMH1FUp1Gw
NWKfiOm5Biy/lUFpCDRuS46GVwpgL3GYkXAcZv8b7lvStXzkZQRXfT/HxrlS0f5pbXafu5Rllx9z
69iiSqv4gT0TvTNqPW6nhhwJos5yMm2pBrTkz6NXx5Bf1DPt8h9N6Fu03ay5zPEYmu/jsCovpNLi
foABPeEuStLwNg/3syQZ/LyQJue6jbDaE9VR0kY8Iygav3KpUXn/KdkMJuGzavJ0Y7v1rdx/psPx
q+v66XVRBPEDvg008fiPf51uOH98QHGYLmBei/7ysX8V7QLDoNpJ+hid1lgN7uTTawqbQKrurri3
jxNp4dWzq8aq7Inyu/sr4slyi6S/jnLb+edi9HwdtN7lW8U8hRIE7EbdTsamAXV+QkuNpq37OqBj
YEwJ8ZlFZop4nsIgxXgElHszDG5+pHoLRFyqq24kWpqJX7cvYKhMmvQ7C3X3zsrK0iTHojFJSAFj
9KLdxc1se47Wi4+hBeMrvnM1a7Kjoo4OrUAuGBVjAh4PA/t/3Zo1GDPptRy6lxUgho0oJCITYmdL
DfazORd4Y0szgw9usilNb7SPAFQtgbu67pt6i2tPZ2gM64otbG00RfsTl77iInw0s+rRDKEpTdDx
3Bwm5E3Ef4hYoTqRE51EeNQ4AqPe3Yi5ZPJq9I9G5Jq2zCd9KMc7C+XmaVbyHRQC6TsEpD1XUHk5
Cf7ymQN/iw2MXPRc+ZZduEXlRBDT69HiK0b45bviiXzabEL5Ru9uhdXn2vHt3WEUUxPCzwR9llxA
rWbJtLqbvHu51a0arF+xGMgzdsyG8mfRpVclwSPuiKYFCzfCgbRErOCXCPlk058xEJMXqvOZUvyB
de00CMwWgpb4TOV+hTMzOlaHGEWUm5Ip+roDGPZymxTwjnb7tvKAWiYuEi26/CfMaq+zF9gZN/xB
lfpyaIIaIxlagrHRpZXM4r1kTXy3tcknsGaExYvdqFmGdjaAyM+tbFGitnTE1RE5+UZdfvfLpxOq
OvAk+RKfGEfts7SPjN3s2gmpUH1tNU9ts+HGotrIuwPgUEcLPGtSLG5VK/GQZf5moevJ2FEmJCJw
l1iYuTQdjk1fS8k72GTgq34TXAXdyiwNBFMFOGdiLVvqYBdgnsYpgGrYxen66I9WneaCt+WoPG6L
m8IayUGgXSBQMSe2K+yvzp423FKS3vWz3/PK3G16HeIxf+dchoRK/YNCPjS/VRh1UYDj24ne1nbl
Oiystp7y323K8L4fhRZb/9AXr8IqNWxX/oBJMd+Yt0XVci63aiGUO8hZvVOX+yyQmd0CCOxukLR7
AO/tdDSIpTfgdsN0nHNjmvaK/M67WOxDtYg6rkCgXift0ql/ExVlivM1kxWEhPJQ79iMHTNLL5tc
Lkj4nV7WTnI0N0Z5PFOr+PCcYSCoge2qP8HhvxTCaCc2ZhJ2ssT3WlKdz2sO+5ShgJYDlPPHl3oU
lXHKuNEqZRPMO1Z+y5zr6p4l+U4HipD60BzOM+wnS+FLNH2zzsa0vSkQfUrIRH/Ur6w7/bkDScQJ
5+P+Y6R/B2oRaQeLBK7rmOZ0lpPZr9IbOVGSQVOdpfD7vmrdGL/EY147OxVuV9ylhtd/5kowUdNz
7BwcBZ1INRKB0OzsYjeCu6YrgwHSNFav3dzufxMKI0TWf/cJUi6VbxuPRmobgi72Y0D1hq5luGKx
ArP/19Hs4+wb/ax8v2ErpUwts47ceNRUqYdw0PT1GeNgHiB1mENZ9G++G/MkVNRheYeqShK3Yy/d
pSqNjlptwNU/DUrNpsZ7lSOci44RknqTa4PLtDouT3L5tLEHMHq4J0BQ2uhtFG5BDCEO8DeTNZVl
HNyn/wSJi8FlPnF9eMQHWoZzn8uL5BEX8SbOnuoyl2tjB3xfAIfIe9jT/Z3U9V+fQuc3Qla0gETL
H40YIB0qHTGMLCVKm7oFYNMsFrwvijkk3UbO3ww+WMmyQ4AZbUANIBeggHzwaOfKpHDwgPPKvr+8
hXScACrEZIZVmwXnCIide0fEjOcyJdLoWpcyDsNKzLGUtBPd3UIrQ9LrVfdW0amcSNUYzjApdugZ
gfDDNOZGyLjutJMxnhRUNGjeUSu2l2Zj8FqFobXpa8dR8u4vbVA4mTMs3Yn1Gzc/v/Ed80Bjfgnw
8JM/7zR8zoaUqmNvVHnbzKCFViq7KkvQIzqBICT2PfDiSQXVayqh3/KT8Jk6UTLYSV3hSb0K3H55
4/UQbYQKIA+SB0EhmZWbY2idnPPxDn+6T9KyYcbPAP/27QdNTZ2ebv9Ske0qIfijTyugN9+5InlF
lWE281353J0CP3UfxpOhgMbXWMMfHf5r09cNyu4elfnEso1ivrsy15hWHS9fDxy0Q+KUK4yE/k4M
Vk7B+8XrjgMwRaebVpeXz+vSKadyPgC/Q0gbs6WmtVzF2/X7ZPqYhV9JJie+inmKdg1ggiuOQ6Aa
dCwSTfE96ejSzpFHENmR6PWuEnRsRV9Ihpn1fj8HkzMq9FOtiySjwT2v8udxoGo2Cm+tP0HxQBYw
WcRhucnWXnSNg3t/TBZcKT/szOr9g8FgeyRVmeeYSUgBzlh8zM7UQYavvX0mtk0I0S18aXR+TiQI
PTi5kZ0ejkQXi9X6567qFcDmbYX7Y+NigFQTIj3tCQ578lIZi7qlDNoHwSGnxTjXxoOtQFkmM9D0
Lljvk/TYvKWNH2/LCDRqC2jITbL3DEvv5gspeAeAeKV8M5b6wBORThZbjieqkuWyrVRinMRY3j+2
VO8S5JWnEwZk8Doven+6PNUsqglhTa2KRJyNye11vUESteavVGxZvTOScQ6sguCuk2QjEKlyx6Fb
DrPxDdc2EL2urn1Dqn5EPkVKL6As2L59MvjWechYt6fJFYtNDktVTpksAnZ4hXfQV9jncGi2I3tM
FR4LjSlXEPj1bKm6jj5EesYocHWMg+6if4xFQq37ntASJpaSFuRjcMlABOZlN/rABCmYB8rp6bBp
7XK1puW7bIMdoRjJrYWEo3xHByXVF3ceGKWiOazw77ivX8qsuUKoc7KMSOuTghZ/e50SWt8MuL+U
kl+0ABjQSuxnunjMGjxMikTayNm/HNhiscaP4mTZLy/yZ49rloHUAco4foSH5H7RGXXOh0+jebF7
Gdv1dxoo3w3qdcqNqK9Uw2toB2f0FpWpB9apn7Y32nySiHc45SFb4tCId0X2Vd21KN/6AwoqwkNj
000cwRxUsTb41v+eIR/BwCkgbIKOIxjeoO0nNwzzdI4BY/elAPudIFzw5Sd4ansqHMiuzTFinLDd
ODzi/PGz6Qem4B/dVaqZqSGl3ItQ6bvq4qGOIn4SnYWVwYIKuOpHGuZRVnoV+7hCtj8yHcwy5pBl
qTUlSMOlxmCYbOa1Xbm5NWlmPkUv3jPwX+BeBNzCnH00yf/QpbZOehe7PYs2G59NOHkaSIvASb3f
iW6wg3UveNYzznvV8XnUlkq3Dy7xfqqILZ9A+K926+Zjn20e6fib/+57rfMlnOq/n5eCZ7FurFQ0
YIJI4enS5lpHiRfrOegu8YF5sueGKRKRceqWTDwIAt3u+FAJh0xqZOwMLe0VoFDoUNHMm59X3iqE
qCNszMwekZS7UVzooORCtWBElKs/z281FSgzFsnfwYLqVqCNnLkm+PMvZV0XHTLJm9p7KkjE4iCs
PBazAgitWWgjJbt9bUdIewLwEXKH/S+ksDZQEKbiv29XbQLqRd98bfkY0RYfzhZlsHiFx4eIqaVc
o5OP9xNlNDz6W1WjGniE3opVCZ3IGJ8GA18G7TtlGLRmgNBdjo/9I13FffMUINV5u8O0zmmjmMaD
DSeJOui796TBz25KnaTcKAmRn/sHI7EOISONoxtyYwMCMe57so3IT97TEPEFhcVEDPWTd/HYvpW4
lXDgFLMSX3KmXFdymI1nAguXqKvZOy3As5+dUY386p/XKnGWe09DNS2N0cKh4wZCgsHm3Csl3WjL
xBj0CKjhABqKGIJk1pp/Id8bb/kre4Vt6FU/NbDGDo/lsXpfjnPvjPDvHj1fLDTfojhu2cAlZzeY
82yoBCR74ZAJaZofxsl6ycjZvJD4q7hXE0dQuZiorD/7Ui/X6sGGpFmUY4QxINxc+y1BPNNmE/31
IbV8m+0immVEUX2PnZqCX8CTuBbvdK3BHMHLsDiz3s8GvSr7PZMwR2SawYR3MF/cIMe/3HrS6Tg2
tTl+7F8z+Fca9762uc517T0n9aP44bQ4x5O21mi3mqZCfZA4je+t1eDRIEZVztNOLZKNER8hYJOz
/Xx8SIv+SkvIbWXbWmoJ5Gfjk+q2/kil2IH0kXG2HH+4+5jAMOH23a5py8OvkusJVCVgvQqwu1/h
4ANzxenLg/EhMvr/z6un+kJzzklB2mui/8Q4ONJvQ4p9pEZuWUurfx2GZzCMlpK3RKNUnyJRUO5A
5gszfYynGw1GH4pFvVqUwsCsTii2kTG2zHLIrBG0yT23Ba+5xJwQOD5Ox6Vfi1foCgbMBeiVihVm
s2VJB5dBxJt36TaK3gMjlVFohIhu4zr4Ftbj+26MzcyHLrRBMwZpXbE04tReHQs4sIgb7f/dCPML
0HgPx4pAdel1Zyy5+Qx0wi37isrXzlXnDSvN//9ZcSHZN6SC08jeDGgFLxfFmh7/d8ia3nEoKFEy
xCiWeBGQFGdzKpyVlWQpjvAUCDzRoZ0D8z7Mzy83HY55dEN8Y0ieHT3Ry/QDq+3ma9wCJpEVVDMs
1RzgPVacCjLSbVIsQwyVDtpth5tUQNrfCFDjcnhPi+T+G0YIBMRCdhJciBSmDMiQGqGWA8RkzA1I
Wr4rKhZMAUUs3xp49E/SqWrV0irU/wuIK5LIWC0PyxMlfn0zEpR+pczf0Uh9AemeTdS4qUgcHDSZ
0rGbLse7yIgQtxbvwNsT9mIu2lUhV4j3E3L9P/uX4meazl9/7SkHZUrfZqbQeeCLylglf7XcHorq
KWTW2jJ4kLakUozBPBhkNwTPqCw4dNP+dXGv3mQ2Rnk6EsCMj8U3TwtaOdKwZPWDs9TGybSc5Ezf
pw7e4vdue+eH34rUF+QrnTmqIEeHh2Y/NE+2RPJKa+DAGQ+tdevLERI9L3bQGU9m+urjR9QULPvR
Ynj8MWa8Rj06pAUUZ/ngYp4zO8b32m8I7qkj3UTt8x30JcaiX6pFARDesrS3UdvS5PaMKBXBNs/l
BJqWe0QNm/cuckfL7HRy/O2mVnXi50BPiujDCWQyVLaiFuVr/3IaCc+v9a9A+eODTLUdTTX6VY3J
TjwKcNJnSMlXV9bLDg7Af7+G1rHgU3UMqnfh0GwYqq1ItlGBpRVKRKH5Zxv6maoMNMe53Qgpj9yR
J+rW3g0P4cH9gqxq3GrPKkDdjKvES69akqrXtYlGzhZatX64OecWqoar5yXIZc/IHz4T5PierVoq
DTt4g7zu0RlmkuQyJr4jRPHfVjpOzcIWyxvO+JFe1KNQOFHHOOkmvevqIxhsCMdGTotBdundDIxu
HaGAsWCHAsVr/Knfs1B+0Q1RBvTBU98W/h/c136MmS69GzlwNugHgjF0ZZ6BmDuZeaWdKcJyYKsm
+lPU/B1NfZ2s5IEg1KZup8aXfEoeXzJrAY5jWZcx/TYgPPwulhzAiC3rTnfXr5KnTU+Z6ELCNdDQ
ODU8UGCwKOtbkz6L9mF+kkhIU0dGvamumWMsLIcHK7m8JJEbJZ8UwAEAhQhkhIQzk94zGw8wWQmA
7W+Q0bBclwISte9n7URdAYFC+5Up0i3eazwX+00jg/sLt9UAkLfhMMvStzDHBy++gMOwnCB8Nl98
DxJdpSM8S8snZbOdHSOUjfwG6lzeQEGx4uDXrIZWcqIm4aTSymRJRE773dtaGEEFWvxV9nBTeHal
sZ47vvSJzUklf5zoKcqWtB6QGTOj6KN6qlXTzWX6jzgED0VN0aLA5Y7IR9TJcDt28zc5N9GKEEfb
GtOiNDDKfouJPd0SdItLbW1VMwYCeTy2FjMLcP85E3Ju3BUX5k1Z/7Og2JZQ7k254KFwXImjH5f7
SAfcF31P25hBXd7mDDCiU4jygrGpS3VVAgj2FRhFhGQNi3s1bjt8fIG5fudFKceN0hTa0bjHMgjL
sqX9vxR37XEKLd3+y+aAHJ66nSIVSjG+PyoXZgHcL3gQt8KzK7+aAOYTXvuS7tnXgas83u2Af8r7
Lt7NHDu7Jb9zSSEkK3+K7+qhtQoTIQyX2rqwkU4Mf3mkvr3aotzBarnjYQx6AQA7wy8UUS+ycU0k
HFUxRSCo3LCwrAd4E7/TangAC/sLINKSUWK6TKRmT9mmQW9Tpm04a3O22QO02IZY0Qo6CTLZMbtW
HFe1Ud4QxHyvl6lVRGf0HBH96+FLG08cZs1zhcn4O+OSw0cz9ERCA1F3w/SdyvqB3zLDx8Ozr7O3
ruS7jxoCabK8AsH13/9meunMeGWfjcLD4hZgQN2vkzH9cvWFsMVWtMmirtlvLS4hQxAoxKfje4jY
Ygq0JMLVjMSzc+eswcvPHTJ0rqHPTsz7d52sDjMn1rLmn+AXO/BLitPvkAaIlspxzjvA800fzuKq
YhLw6Oqm4QpLW7Gzu+6ALh7khpfndgGgpxsXlITp3ziP4xUlaDp61FWt/TDL+LTMPaU4WGQQCaHf
NOfiqyc4Y02J02QsCUFg2X08YdWIDKzaAn/EJJ867YeEPAeRxolEZ5ARhBNKKbTZYVDOlXIUq7AR
UiAbkV7DAZ+/f4+btlfe99R84sf6yu8Oe0hEEtRckBw1r8wE1VibOHW4mjhzx0Z22gSrIdSI7vHB
CHyh3g7GyGJNmBlSWzcSGAchBX7lgerlDoFAJ56schNctzH2d4OObd0GMbFwR2vvQfY4pCxALoCf
1sPcHAz877gxyOzIWJzh0iOJjgoaDdGOu2f6jBgKguO06qwPu1u5TtF9Yg7pC6TUq/ix0t6EC4sc
12jFHOzqxx8GQ60LBkaZllZBjcxPIoMOcL1rb4TfM+C0h+cDvZSqGGE2yiGmAtrcBtf8DU34v4Fe
8BLS6ScyZb7l+qU31n/MQGCioKlezQB/uDY7zSmt3eiucVt0WPUvmqXq4i0CvfJ8BxcaT6CkaM3W
LpUGVbEroO0Shu46TrwW9LOmG+URzMOtQkoP86Qm1QiHMmXomGIq+JpKBMcyPAARE2rtMLdbQ5LS
FmQKnBmVZZh1zUb75jPj6qpauFhzcILoFrRh/UZKMSD+51nFEMf5aPpWXmMfCtEZdADHyn19jI4N
+s5d98aYrzF9xYKLS3czN3U2juSRrvUD1ULRTjE17Yy7LhDqMmCYlXkF9nwScYnz04arOEppdTBl
N2DDtcoSuqY61QwTuVFAlFxkHxFYEmUbLANkkZVPUKxlbhtfCldh8mT4oltxzpDyB8Zw9XXkMgEV
eHo7uN6zFKvj3UBIzxoyqP9mF7moip1o7iFD4lip2gFXKp7THYHSRICcmbebA29bPPlLKBzzSQWw
Y8U6BxdGRAd1A6EtPG9Bzw7koShXcPV2CWOAYFHLWLoApkZ5JfNzGo8dpOI3Y7e8mUo4vGAyfLcG
ErYHIlZWFMwJoIQ0QBZkrk7E2deY6fZKt85qJfR5VRa4EihfEZUlVrrcGkuzguzZvHSI51xerGOA
rKTy0hyrX11g4UfXWidOaIdgBMlIknG//SLvcqJ/iREQ7kp0Sg5EYsHftrby6kW0mPjYH5Yphylx
6UUb0ZMM3d3UGmW6S0E7u/RDB8Ao3LXM21wAGqJY7rBT/57OVuvNXQfmzZDPBlh2ICWACpPTA8l5
vbOaoDxnVQbwCgQgClWQOcAKaFR9f7VmkFUuVYg1eyRQShiALXqLlCCOqxNUC/to9hJIMia3wG1Z
N7vx+Y+Qe4qj9MYxetgHtB21v0Gh58NWtVT2XFRQCKfjXmnHhU7ysaciAmVYFIJxw38xh93eAYy8
Uq1BBWSzW6gu90JZgbnVVRU6IWvRB4xWs10Y0FYILhkUgNvZPQYhqFXGyKwEDJLqROX8tWuBF5Ng
5JfLUMJl+p3reHVk4ZKPKH17VpPX+KL1EzxQdIxAlXpCbCUopNq6WmH4p/6ZQ7vFtUAKNrdFSeqD
e6tX1KfvmWKSgoZTXxPwt++FU9fOIONS4D2e6UNgzXoN+zRKqYaydTqvAEFyT9aDS5gULfAu4Fpw
BKQlJ1/xf+Cle4ccuoUMpARIdsYvDMcsVxj7nIIfqkCkO3wtWOg0U1semI8PCvEZz2f8zv7X4hVs
Jg/3FXwG2jc70tlMRfqU2r12uHqGHaZdMn6Pxce830CK0QfoQXTjcI115fO2bDNPUYVe10JOMPuP
seU19NVTt32OJgA6/1TnQoA78hZUNNOvAy8Ui05LYScLI1r3JtslwosHXKXvvQNtblNPXmrrgITQ
8xYcVv1RuwwJMfEbkMzgcJokwfefRL/RhnTewEudlv3zaFzQ5uxrovFmSdHKn2NJg9bOO4vdPRRo
UIE4ncKrOwnucGU1BqEBMnF3RM+4djpHM6iNBf7/hF+ej7UQS2sxxBZP8cQHnPxq63+tjQ/0k/Zj
mQFnJFmGo0MEMIOxrxtBLXjsaX6PxAN94m1CIYo+X0WWcz1seD+BB2yJCYF47hZI7Rgv6r0eKMsz
Zs5B/NsAemZdCU19YgbtSEmTVWhd4RJD7FGmtwX+t9U0rFzzJLPsMFJxsq2TBAFo/3iIPQqbxGOd
HtY94PQB9Z9ragQFQ1fIIJ98Py50PYG6KLVhDNXLOWQZ+GV5GKWFWlfwq1BO/hYLQx1BNiCFVpr6
OMLsi7sX8v5mR2qOfIHPguOaV53TV5MFTkBZk9k7+ty3Za+t1bpT0Q3oQr4exQ+KWitNoLApe7rd
C+S0stzPK5+D63LpHwoHvuUioKTIzRtY9Pk1gCgxd6geLNiVVqZ/VbPEvo+/YmeedLkYsW14P96d
THzN6W/EZhFCLftjOz9J8c8FC4rBLq/3cd2eQ4sIhOktquFKB4oamLPb7naBIF3JPFJqX4jCHVkV
MWnsM+hQCMTp7O3qi2F+i+MoTHUJW2uTC76A+21izzZWJP6jAsZUUvxsVdsSiZQpvSLSSnT1GWwc
DOS/PiHgga1ULFfO+C2FKLAB7hrB2HwsjTclFGAHoiMo+3OXybpKgAbO+7vvBfp2MwAreHhsigl8
KLtL1bx9tPogTU0UihZ595GHbeO1M1mPL0iFUnC09cZQEtR9hll3BeQUQXTA8sarNeBPjFLdavGy
xXCmyGU5LaICaPB5+VhbPCnLg1hTnKeycHCZN4Mws63X4jG1T6SaU9gQ3zN1fkyLTQ8LlCBfpzi5
I3ip/9CyWMEz7giCvmQgsK5sZ9xF0n9DAlqCplq6j0tM9HTLF1BB23wnAmUtYeljSWlQv8SpdXCR
PtyNmM4rWL3S2ZRfVNPgyuPKO7s8htSWGRpm4ZXHnXbqWvVFzDsBTALtizOR/2GZqXjHyS/l5CKO
jyOLBcHo7QBpKrD1zV/KUQTZBVAwBb9o2MkVHSYPxEJ47vnofsDvzs67nMVw/spppCqnLzd3+5kQ
Hw6v4sm2tVLhCTaB8n1YfJppgl131TGKHeN4nt//DdSMb8kZz+JcpJLWwyWXADn1hHSBb5k0mQLG
SC55UMeeaqIkqhqRlHSlQ9gqZzTvvkSmHzCc/hoV1GA5Ww+cz8m247eObi5MX7sehabLqrEgfQ3k
0jt2T4/Ze8Hg3cID+JxmQfysaYLbP0Qz96qXyXE3Cl5LpMrazJopLg9tJagokDvDsPUiUxBCKiHA
HEmvxy6EZqAbrsbXn8sh9qeYSGmdKiYguvZH0ieM2qcZ6xyItS6/btqT0C2kAM00G7goDyOtRLS/
9vF8Rthz2mrA8zSI64hNow9IABbPOhfvxtUThzUkD4/sTEuFC/W43K5g9i+eS4rL9HJ6tJeOPGVW
gnDhE6Q4X5cPh5Bz00aq7nS/wdldltEXUj3w6mVJewNm96L9Ex6cjV4DMWoP8W82Y1nWOXWoyljs
6QmEfjNp+TBoQa7LhJ5d/i6NAsFn//oRBYXc1ff7zwNJ3BA3LI5JmvgPeiujzrRRJvfqDpppx78T
p2p6mreiFfZuaa7VaNYZpTOl2gmgIhSRuw4FZsXAbF3OPbg1UeFLHgL8K/SZ3CREj0QIMQTnA0/E
0Hd+xnSIds55zXBVl+Af/QLwudNtKQojXTWqH2M5vc9wRJcvLCm3Zqfyn4naOZ4cqLcWZNQnwtQ7
UrL2IDtWHWeV0X0EyBdw6FwSWtKQQ+H5O+Mszv9hQBFV5DHGRW555ijT7sugZllFMuO/rK8ZJw3c
VyZLiOMmnM+mG38GuRgjcpgiSz8ASRBjMXxIvADoOq1j/3s0HvxvRJ5zC7nkjZeVkMkUDkmJGK80
st+T+pAtIKFamDoGM4zpQWh64M6vANWvBiY8TZbio5wxz0Wr8ln+f6ip3+/d/1xm0kOLo11dzWmb
6mQ2lol3UbTe9QNRi2qZh87OOyONnMdh8ANBvgwEiTg6IxAS3aNTSSxDeMlxRnf0qp/id5iXLHiD
YUaLHbbfVzu5eiklTTWGyCdhv1gD480txMmogWkIiCnpQJ5NyTeShuxqv4NiL9NbFGnUjTv6Fm2v
ZNlrN4R0+0Pr3aJjcqj191njskW2cT1bWLN75ByU5yEBQ0ZyFp1uvRQxwH8nOVwhmk3Ypu2xsvyK
soohbW/Olt7MxLfQpXRgwYQ/YXkSkOdTxVXrPaRDQsM2hUp16HdgCBtxYnaNV/PSs1CjzLKUtiMz
LNtYK/3xp+fCZuKeb+9ODHHfE1PFRBa/7C3K4kGOvFt/w/l1nYM4s3JNNGJiTi58fFrEMRW7y/mO
gcLk+RWIbqhjHtb2SMbPqFEsX4ZzuxJnTk6EGi/ciu5qCBIpmeqD/iTXTSatUU4KxbSrx09h1/IT
oSk4yj9VHiDbEnoauZvD5vkUUSxzgqmO24BO13Fbsua0uKTQIbKfWPLRq68AUs2JFruB5h4E3rdw
MZ77+lU2KfxejOkyDDLPKHK4dA9mGwehOjyp+//rYSCFr3YIeWvC7fyAc2sf6iBh1Xd8Ef1DyQaW
ESmGbwVaUZgkpn++1Pbd2BN4IXxDBB2FwbO54ntYWp+UfkgT/mIglgxY3Znwo8q2RjWNW21IDGPw
5e4OGkxtRC6kvcXae1xz7lGhwLvgOby7i3prhuDJnLpPcX9Zxoqv++pjfz0pEY2it57FkxuN1Ixa
93a6v0Rq7RucPMoHYvuD/klakalmR9052UOdm8Hfp099F09zMdUOGkAIYtgOTDkCTkYuuaror3aw
ALh7uGC7BXrJtW2Cz//Z2yoFaNsUcLQHfHwrlANakA0Ga48CilMtcEg0HqNsavffMRD68eCefN1T
XIuiZZPyv71ViSjDd/KyT397vn+/N9Hq7D85QDYEnprjQvtB1IrpXx4bvW6KWUgK7LnXycLWMbEr
5vA5zW6eVEI8Agfo0uQ+kur8+GTyJ0V10VJeQYa5h9JCkAqBA95hLQpyTrOS60eGXyvfKcUH7rQk
e48HGZEmqPGrQv0eaOo4GkFtf4YDsyKyfARAGI0hP6e2zLPFEnJD7CQ7itQ3n7WVML4ew83kCdJ+
tWfWOLGNhWipayV/EW+89iUUST0dMwZK9c3GFHK++2XFRB2zw8Dc+6adrmI97utxfe3FLDlmQsNf
aLEnqnGs61QfXprzihEMG8NYIGHoTu/+r5i3w3pwnw4wcjPw33Vofma6HsJlcWN8F1AxiokNjPn+
zXYk9ovfVnCTLdzsgxvdQyJg5iosvrsIlnzB9H+qwXsKuEScEvTvvh3vY6pVmgIIMWzPxgYhdNel
trQkf1N5nElzr2jzgv9vrDTUH16uEDm05VdCWvR8/W+qBcJlot09c/Cvl7NR8zVRKKluO+UNJ42Y
zkFtaj3xSx4pRFiBRaLYLk5lgUeMmVjx6wf+YHXNl4Wzs/RXPx6q5EYZVn1rod7uWiH8i+NaINqa
LIgswbDWrIMkdvTEJiEFucHDpGOqaTRg3DbFADrXFffxDPA2RrtyXpe06iw88TsNfFlvktjYA4JI
0Xtd2KmEo5DSsZ845nDlStUTQF913fSUZnNQuyj9IjwihW/BENSipwj7a7yYP5b5adRm5oP0D/Nz
4K+Mb2GTcEDzu7nZN1lo6oqVZ8S+1I4h4DKYcWRxkunsta2UQcwlJMUAzDsGVOoqgxwCGeeWa271
IwwS45MyjhYU0VFfVpRUB84U5qsUGIMfgNCiq1KFASWKDEk/L13zwp+tmHBrX8/Rf3SLxc53pe0z
e+b8tvb9Wg0BFphtmnkpXRVV418OuXv4BI99PTMXGOmjVy2csrf6WJhtP9kbH7z7xN8txYeI4Yru
GK1VG3CEMSgm6PagnlpFGGCqEQ1CIGK5TSOmoTmOMUzE37WHEy+VlvOMGLPm0xCbEb9GN3clfLYx
ILH/pEWNTIcbH9GYO4WXbLHFNHP2Nk2aJkSbiZdnttYk3Y9T/orjISQjfkJS+a1GAoPoy0rS8L4C
8ZYBDv/Y6DdomIoInFUd6Rkn2E2UPvcpZCSsaeeqUOA/wC0VpFeJXPbH51U43Bf9C8ZNmQUyXeMD
8ktl7TKi0w68feJK16ahHZNBjx0sbdiCMpbRE/VVig5l6+DC5QbubgAt7QfJ+gSwSBA8M271Uju+
l9MgjuGRWeyeEPQCJScDH4tw9+reHKqx63ZsLx6rY97cfeCSTOH2ZOxl9YysK9VIpoLYwgH7GNai
E7aQfp9BPynEC8wXZd6MfZqqmIp2VEnMAsnuv7sEhU7Z3rfY/GOFaz6hSaz292v3LmRs5i5ZvoMl
u7cm1rJGYkYWBXvvuImQ/L4b6Czr5zGgXy7l4a4ros1c/ZLmQ5sH62wFW1fkUMzxA4TU6c/tnthA
O0wyHhzw333i9GrvLGy+oJmVVExIamb1+Vqio9tm1m+UGtqWw32/SwFzUSYb5O8Fg2bMbayjOpee
95MrJ4WTwZKOOIyicOGZkU75/Zk3OhKyYbN0b1K1mnLwOF1NegI6iEBwI3DQILhP11XwftiLGyKJ
hgxIJzJu+cc1Zc5QvkrV/gESNGDsQ1RX4wjnTQ03kCxg4YRHlTLbblc7VzMgseZciGKi3epbMIBl
x2FkjmQx/rr0jsvD2agHcypw8WqPE/ixfQ+twNyBeGUZh0BVlBSvOt1F6W3rzKO+p510mqEadZZA
LTSvxpPsU0q4Vff9Zjz1HtYLZ7JSpujRW2biZ1V0a12ogXNJGQONkOViUgvoEJDu9L9I8Rzjr9C3
+KuNSaQpnXZb5iSv9d6J5i6a5tPgEY7nkJGHzL8tARX4LSaRRoTCQ3kCeQKaly+7T1XljqLqZF3t
J6wNMsOFErERMSzjthkjNEFLzHHROvq39K7he9i+Z7U5BBt47WrdBufQIlbZznnanJQE4mVobRUY
KQA6xoGom4zu96fn198rd/erw9dZPK8hMexd5RVLJNPymv1dU0LWJHx7Gh0FtbT2NARSm622gpJd
N5XHXL+opIgkWDLC5DtUbv7F17/jtGfOQhJNubvPqsGhc3AgDEP7suGQjQSP+NxpqW5t0jLRn1gy
hBnAiWqEUKm07u4cHGnqcskdXuE53CzeQsNvscO6z8Df7V/NavH1ll/6yt9RlSOTthn/qb23fCH2
dubkoFI7UVOauymT6gwsjMOtGSLHLfFzNe6BkDTcF+65pKGIBkCsDcoM1btx64js8QxJ3Jxq6b7H
EyjeyHvzTJYBR/XRPyrNwGJjzhpOM6W2kDdOcf7UL1b+FtvkvK+a4AXk0IPlVvxZyC3/xryASOKk
hNOtTWhHOc0gRNXwhS9QMVyYx8LT4kfE0SpEc6d4P7LPFm0jMc0IScSfUFMyS7sF8jKWOJrl2U9Z
V2kaejzGLMEfY4KWKJCBGZh4itIt6hW3UL0QotNdmLSLUGf0nQtIMpgqlBw9EzQ9aNmP7PqbtOy4
o8CiK0v9kkl4abCadHDIaMhRSjPsohsgu8rATWWOSA7gsUJNTR+GfMIasHdIlWhhPMVsXXDJzWTJ
jQaEg4I3IS4Axy+pPJsQ+mp+klECqIz5x1qTd9mfesMHI71EZ+2tJX7r5aZfJUpHYGrC8saIOKBj
kgkmDonRlEnT/avBtKz6jB7vDgaN0080gRsoDuYW/BTcsArhsvqqSEzypv3DUH1tqF3Hs9JoXNgl
BmGSRLdaF/z351/KpIoiCempsvGt/4U39im1Z6yyzTij9m6MIi9iigyAM+vMK2+FEQ3jYc0bw4iw
cs4gJcQf4o5jp12KnaP0eHkZbpBl4KwuXcdy6p5u0Luz5vF3G5xjA6h8Mhrgs4/FGI5s9n3XQFV2
rXNWvzdfauiKDUoXUZ4+0LmRyBAzAkWfDT5nO3fTPiHdyPGKt0qcNQBQmNjOvlEE1MYyekBOTNOc
hh6vl03v/hvGeMGiHvUIRzVKVtyFjcBRng9ohdX9Z6zk5BR+YUPyIiNDURn5lUeVYmiFcI5VWFpb
4so/4ZwKgkA37z6TtQ5XjbTvKtMuobDax5cupOxXPg0b8RgcxLg2FYiVCUuVWz/kVd8So/w1auwF
LnEE2IrDvoL/SD5wtu8s04S+TMFLfSz3XoK036qJwvnqw5YaoZoosvbun/nk2p+rYi/mVD7i1j72
Vo0qxLCWf59V2Fe3vFgR6MFnR1B5wTP7s21kAadTnDMLBkiBMf7Xcx3K7jqyPXJca+1Une/r7CxI
x7oG9mQ0HRZIRAAN9J4SKVRBY51P6dYGZybMDobrWMVW6joLLuHR9RXJ7cHiSaziMGlwwok8159C
NGJr2WNQD8wdLR1GlS1uhqWI9+Dajy5rQfBSMnFeEiJpsvMdJw23Hvo+X0xDa5gx2BsqqVlfEnnR
E4zgs4oGVDHHXOeKP4bfpwbcHy2Cu2xytgX7LQTZ3m3JCHNHr325PP53zsAbor2usEhLGlbbrv8I
LEeg6FplTy+djUl+qMVicQAjVz/zq4zomQI3v01SUitQyheNQvo3Pj2XeHQjLJaNUuFoX/gSrc5N
ftyJF1izo3RnUk63fV0rRNcAaoIkuvixrVs0+8mjHVyJTHSdYU2SFEvmP9LpgKPH0wVqbLxn2aIL
5zCXka/lYZIHsc+y6ObBx2JSAGTXkIIpEhSDlLE7q9+WzHrC8bySI50OxCpWS7+C8NBr7iEid6Bo
y1LwO3LCsiGFNMUEKu0sgQWJDP0f5S0xCMfZXAqkkqlKi5zq970wDWaWMnfiQQINRatQr/p/oXUQ
1K20NY0id8/ku/t6rQv4nzDpMs1aO20WIyb11gFWQ6kBVSG8YoySQLOYpF0o1GziS13Ro8tk9Qv2
j7FZDNCK055lGmxAJrxPFKX2mp1WOObarJtiYDBHl9YQhNNZfhKR58a+dPnW+kNp4jGYcAmHwv3w
3xdWsxRrP620+TqiUlgdPBnK2OjBM/3CKb1BYvk9wmAVHXzeocVODVa84QlUnbvulIOuPNyIP9OG
nXhV98A+m5kRe7dvLMUOcmSHdZlX272WuVliBXPrLlal7HOSpRpKZ/W55e2+RwhwQs+A/Yjmfa+I
gkq/KtVeKoTRypmVhrPZ8es7Yx0DqBgBhySiKw62lKFGx3Ktf8zdT35lGYHb7mPO14VEpoH13yLu
lVKnpRH9OVdoPO2SJmHqltJw8vWH+sohvHFthH0fqYJlqwvdttvtsdDolzWJp3SmN/Y4CHSFeI53
oboMyB7vtvY35P+cEFHuk1Npq0atbojbhKN1AGrNr+FTjvG7HqrSdpLd8GmQQovEwsTWfJRqJw4g
30QPmdNgOvJ1BWMboLiDlkwgJFLyB+/33PSycic9jLZb2HhWGyYnpbLoEadM0JBlkLcGFgTMKHgK
i0LhZ6fpIntx9A9mjW4GCwz2G0nOkgtQUykpCUKNs8g6ofHSO90q0hRsqi26JHow98jwKeCyjYcT
2aeaNoztdIWndwrW4Om8HQ7b6A6EA8XL90JnwVNiIxdo/mWl+FumMsKudJMam7JY6lYqM6RAqRLu
/hXJJ8cwLQ+MU8Y/ce02s84QELn/Mjyb6vAlfRJbLWkxHbPE2WHdJAKiug167p8UO2AgmYKCYq4K
X3fxPSsBnc2h4xbtPu1zL+cQFOnyUJ4vaOfTmELGD3cqnce4Xok59Dkertoy4/TF+rUATHMwf+wM
b4B0r9DscOtucMD8IFrfX6yPh7cFT5YGqUNA0qegmdMX6RjjR5hLj7UBdn6rIkhAyUPfKhbJJusO
1Z+RU/4j5CS29B8dmUX64BMDgtRPsZ5Pin3E9yEcgWxvwRjdClNZ1OjcgEsU1ENNy2XXaUGacief
AhC16o58xaY30C3KJ9TaioijYUQUHQ0g3t9Vo3AtCyKOFlXxDMlCI3ZF0kIstdSMD/AflWPRdmmK
JTGGRDu8utVW812mLjeJU8x8hiIIg89iMXgTdUhXKq7hgoWqO0pHzJmjBsDfXk3T357iIDMdEkJX
/g7cAi2g1mhvzqT3yg24JEY3wAFSNEfT+XyR9uKsOIGRNwVLJITIuaqPCwsaz1BDw3jGAXBCKso4
9pXgGBzFYLXA4znW0KxAwfYmpD0KebHkxfBGh2g0VuSyDBGivdGPW2oA14ziozhVqRdPV1PWbVOh
mwwoJxHwYWsi8rrunZYa/j9FUkkCgpJnTbixuefEmYt8qV7uS/PmHRe/pXiU2/1MJhgxpsIs3cAy
Yv+zAGfmSsDz+J8I0V31PTCmjBZdc0XrSQ8Y2xx8lLiRG+YWAGkTAW68aYxcDEarIn+xDwJMi+lM
IgCvTKm+hG3J/3ZBeKzQFe55Fu7hzgLndnRr07lDFoUQTUfZ7Ja9vPX21ix1kw3JB12AWsL8MZ7w
0t35aEXq5hJWWTGgozs0uaXHZN81bvIMT9BoNTFtPX/JPUnSy4FjPblLsu7TLWWylYmd1VDMB+L2
ONCXo6xzJF+RObdMfxgYOXN+vhAMlknoA7ggN+07RSuFeDXSKzo4TXJYDLqjkDYty6T7xJYcO91f
B3Zmu4ikiL+khXdSmYecxxruLgNhtZY6xyGAxsnCRHjcDDyiITj7gHrA6fCyp1qhXiXIDMN6cYec
fZjJFcS7fRpPeR8cdpl8qvuJuJukNpE/TMaxhtpBRe+0YGGnPl+jCeA2s6w3tT7dhC0UZA+WCqE4
ga72d4ZUUarTx2oo/OO8+EZhCmsm/emlwkKLkt8ECQx8PYbBz3EYDDL9RlhhjQOcaZ1tybnhuU5Z
5fowYTuQhGeXGA55sZvpe3yw5PfNh8ahrXrBz4bJ7quN+gwBfXpiz936ibnsZ9X1oEufYVLVU8qE
j+EJ2UcV3tyNH5leblk+okz0Sy/mfFh1z9XiFQ9B2GeFnN1dSO8hGDr8A/OjYZSumajpO/GpfuyS
MKHzoqPzTSly08wMltt8xLfC1DKIa/8bEAZ1i078YZ7NPoP/rc3bYHgbn+/1zdraDwvkdTkYbpos
8PLInuLgw9qabIPfg6m/wYF9ZdCE1kdsKSTpmf/QCHCLcmmT+5AUMJ8yJv/qcCtnBx4S0F0vEjSR
l0dnCPaG06xU3XcqDIG7MVqx+rIa2RUU/ub/CkiGvB+iz98Tcv9sYNRF46SQUmAAB5gc2HtNzsnJ
5fyyMp/uUv2y9zcxj4neXPpEDm5QmHXEfTlR4w+p2QdFNRUEM1s0SqbrkRi5t/EsU0B+sxbeNH3X
aNt1siGGkWci7l0MOi1Y07trBWQNcDbyXlJBk/eFZqMJ7BaT3SJIt3+F52TS+HogXtahZO+RNTEV
KL9Cg0BFfHsVCLiZzr5WJh9BRTfVFm4l3OpexLqn84Phk6yAotOc7bBVM6vKRHCZCdA6fzMAiuc5
f2I+j7qjERqun5yJlhr957yX4n8fhCIaBPe5iRvX0Gw2FgE8KAi5cgpNkxQ0JzHRBwxkwFvhiglg
KKQmSri5itfLnai9mvXw5mEbjhT4/7Gb5h5gWbJ5i/sdVn2ZLalGHOKoMsoZvd5hd64/ee9MMDEK
8RmwsCsqSI9zYPHVGaXLUEalPrA7EIpieI3Cvi7ywHAsO6AnSwoSRaaqLL4jauMzGwYQFTlWq3Hg
thW73vbS2tH1MDWPuPjTByudDku5NGv+u4U88pof1gkS//05DZmo7eCLf9CbeP1tvd/7pYbIvmwV
TuzbKjj5neI/djBRwvsvA9pB5Zgz7SaiOu5yqDcqYsFtcF3UiVm8cBkXkNBea+Xlc189W6tWIje6
tlqEGuSqj/8EY8ehYV6PO6Kdk0P0gkCbT464yd3FkjdxBnGbiHmw/aL+ott/4MQhMnIlvlDtNQmK
dFsWWuxbnHZ0BChbO0z79ROwbLD7waOSvG0PeWvvdeB8ubFfEhSYCuHuVtnH4yUBvrd3dHeJ6Clk
oYk6KHmyDHzNg8qUrBwk8IaroJ1yg21ZjjECqUj+GNASm6Y0VSt2YeLXN1xF6fCHa2y0/PrEHjRs
9/n8JLd32DnVxRHBRQp4OcpuOWSdE0EIIRTv6jFJsf4WCL82YK7m3HMBKpJvYE8+RibaAgjI08LX
YdaVwBXXyRvmMYndMFN3KN7bO/Fjd7yJvW6dOwwSLjiz0r9mU0CKLsRISU5tfuOY31EU63KuI2mO
KS2QveRpZ+39ch3QRBLCjtgsTGbzj5Ghtb2n9YOM5m6E1cHOD+aFFj3LXO0cxoMZ6OjgqeUhJyJ0
EwK8FkxzlRqItTQysIWYWPEHXyfu3qxXPktm1Cx+hZU4a4NDQKaFHjUavAlSyY/z2Ys6LXgMwv3k
8hyx+KfKfJRSMFLgmfS90P6ktx0w3E+pwnOoD+F5UZRsefO2T0NeUojI2/Ry+OhCHuEGdJkM5gvp
b4rxnlccv4zw1IWL1H6G3iVH1HCwuQU0G2L8pX8/OOzXBGL/VxFS4ODOylcuSgHFiKvuZELbJqAu
i2xvAHpE/yz1P+2yjuXt02Eqs3/DMP2JWOWP4upxGFBbVuTqoVG5Dxfc7Y2hvMFJSw/ZiMM+YZmh
7s1I+nH5Ed7MTHQyzDPMd2yd/a6UiLQHihEwuJbuR+WoEcUSg+QWlBQVosjGPgGNiSBYXrFdoMEJ
QNOnTlWRLsck9iujonEEhO9/L8OoRwPw6kqWi2TvgT3VCNqZ736sQ5JajtgTGRaBnYoG9r7ai8t+
9JkRF5f9Wg8tY8bt5nh99cD22W3yc1mRasXtXcjTrHzekYL+hVMWU62C6X0DGf6+OdDpUEdVGtLa
A98UA3T7eQydpGUKc3C4A0CypK9hXJf+HG6ZXxG0xBiWgcOhb9HFvbW1d/k+bAtejxSd/kGTvhD+
XsZxc/Bp6IMBJXGZsiEMJdqdpFT/CndvH/Sb3dgUvV92hTTRWEcvCHF2dnsSqzh4VT11i+LHuGcp
Obbr9M2YBHUb+raAN2PjqnkhKIgvS74I5W7uKhOd8uw+UNxJkfK1RB6g82CLmCD7KXWwD9Fax30W
i24hZm7YJaM0636jYyQntmxWgz9NFLUCTeN57veWPL0clgLgtK+sK7ZcRp/JDHrFb+5ayRgQKtmx
+7h+uzKe0lrGbcV1/oNfVDee7AjCx6Bd6EguTBfutV625I5N6/PLhiz4tnOA6mk7skzNDRUYmbTV
n/Ege+BzjvfSoKpe64ehTQY000D/TqpqaeFrgeRX9HX5Z3fReNW2aK/mgHk5rF41Ie3gM9MsMYM0
5ti4L8wfbgCnr1I5rZuLGSHA/qLyZCRZwz40P3H7erhflavyJlkF6adjmQ6jiwGhJtBOR1+U9Sde
BUyzlOeVKxx5AiSGIXzNIHccDHalN6lt8Tr6x3EAv/GQ/2+/iB2CKbbJonIJvIL2oK7thH1NMkK4
3T6/dvP0dixXUK7rmWGgWxQt6dkgK+xXxIkI88LcRZazpQ0J928gO6OE1jmexCx5/aCSJnyvKymZ
5TNzWlw6GnJDFgfY4iYsfseUXukb9FT4vQAcZU5FYnagKB7sbrHUG0zoYwAaWXHRN7HAkwB0WqnU
qrXFhRmFBaIQRBzopn21puLTlGuKCFF630dREyeGy9Q9FuBtHcDOdeDNFrqytwkPSTuuKT9CLeNs
qK3p1CdNyaHaykg4RRSWV35ncGqEHrp0oB50ygprkn35QYlwcoTAiqdTZuJ5HYFtqkCiLgE++ORO
2szYyX2aUhpauJL1eLO11xuhsTmuyJGMKmMCx9ik6OfeObLy/sQ204t7SmQbkW/aN0VtbHClzn+4
39TTbJLMToF6nUwKYKRuKNbFXTnHnXFYPsvBrCleJmk13ZeBkGNpTOzj8sEv4xMBtlb8RcZRJ2yC
xNTq5tzhgcqSsx77oRGBOHWcx+KnigOTm1erdmHrnWHOazFsO8sZwoVjTUM7VbFrsck5Fv+v+gLX
j+ARBtjHcXu05kGY2gXlLYfVnPRdylB8UNSU9dyXN69Ct1+1aXmvueFu/OT6g3DDQbSj9MIGJUbd
tMcrLK6KckmGoHLehN+unGXpd5+imHYjfv9iDNylQ/87nv33P2BRWeHgXzokHVrb8ZMtYgGPdbRh
GOcJTULuWx/Bq8X36gVJeFoackZwfT5tO4Ok7Bmkxlq1unryIrLVJhB+tBifH4MuZJNeWwYvU6yN
/7CTBeeavMP9EElPEl/XF2A8ZZRFYgrEn9vjE6gm+YiHwSRyrG9TnY0BHNng9JcVbEVqk1cloZ0U
HWp67fc905xyIpjIqxKpdgLyLIJGzKhHhJ0/HxQnB/0Te7DllMZXpQ8KlBuilqxw6TizNjcXKrtq
QUS16NLkcJg0klfqB6jlM+drDEvHZDEJkgKUWIZq6IHKNIslpqhFbtD9c6NOFQZoyT+vcToVN2Fj
Q4L5x+eH3E/B+QJG9lcndv441hFbW6n57/tjY7ztnfQJFdNpwGFkp++FaIb2LTN/wEvlm4+OHNyW
rn2tdyKIp2Dv3jdFRJpHc1NWHy/TGLtICPM/M/YZby26ElzDIaL7KxUZLbc9eMt+S5ZAYeVnjEwJ
u4RSW0jytFbtpt/r4mpdWFaTyVqxztd3xiY4uDIekPYYzjYeWJesCnzwDl8SW6XBRhvC0GjFq0sS
7LjzC1ZvWhSoxRiSMEjIMSJgDHximRYZQBPCA+wU3xgNuKd4ZVhD37hciHIvka/9ITJdaLz/vGdo
8/dY4g3jY+z7mWhDSx0eSHD8/azCuTu/ocfGKCz48yVad826ztLK77siXHKrlO6SUiZRY34PEbUo
c7iDvMRAM0btzitOQviXd2lfzwf2FymjXqLoLNxZ+WWvkUBnAgRVO0XjjIR0nGxKnN4OIeaMPgDc
41qN6p8wwf/DRWKd4Xg4odfZBMAJewfB+mGqb01QTAewJCQUWG+A7U1G+E56Jz7T3bc8f7z7sMqq
RwjynnvKvfCievOUb8fy2wbDO80KlQwdlzuYTGi/1g0A3vicXuxbdNXSvwlzW3E4CP2+/pwDHSFM
z3vGY0KN3M95ky1o+kgOiMWvyBIOI4Wu/GdiGoYCdZMa/Qb88oI25QP5mObDhjCn+Fa1XOTJihnQ
b/C+10xwPnwdfGVhotfAN4Ngv74XzEiMsCxP+PRuYHck1YHOFen1ysIBPODHsFC8ZBBi2e1AKd2c
JTfyHIOJ12Y857rdhqug/Aw+23KCbSMFpwxCqfoLOA2oByyPcoTucRNPwD1ux/zxj9GDNoUr43ey
z0fJA6R0D+E2rRisvxT7IVczMaoPBYEVJY+OsH9EfKyZuE2DzDDkr/YIffKIOTpbDxJAy2Bx5Swz
C6vGkqcL6KOKbv6xqtM2icj3tIWPgWzVc02ZKEw6VJ9AKuZ8apLsej7ytn0A2BX54fATLL+MQIeS
tJC1CaFybvxpuR04sswrY5j/m/AFLMPWYZjb2vV2JPaCXMhbWn62fKwf+6i1ELipc/JXYo3oH3Ub
/LOHAhhS5Fa5xOhm5qV661qsYHxQCuniUTbe5CkZyFmM5ZEt8vJd0X/SNk2yZu22nj+QIAm71EZw
L5aT2Uh/witgJhr2vOZEmMwCe+srkMV5fKBToWCwNbX63cOAtPrar8HcdE0vCBX5uVqnAJpUxrpU
btHOAJFyXf8KY/bvjwQolmHkjhr8biHaHsg4REm7R8KRfOZUeUldnq2N6/PE3IU8fPMAhDs3iWKv
gakSLsMZd4Yc2E48Q0bWzsPA6No7Fw1HdJ9+UHYLOV4u9ivYoXyqG/06iChvuSlleCaQh4vW+6eb
K+hX7WyUGKpruhbIHir1cN1UX0Tb9dzKpDTu5I895EYySti26LHeikFwPR6KIGidu8vEBqErLUia
AwIReGLPARr0r4fNpyqHjNy7jYfWU8S5Al4RjSKWCQJvf7TcRpZFPqrcO9PwS4ySoj612xNSWxMf
asefbgiti2YpNgUTCx/S52ecJpXhLg+X5F/Q2YhBDK4YFjd8Lt+Ga3q9Qum0Oi3kPHMjAqUz1oGx
MhQCHGrqTSNUxPP1ME4lvEp/v8yCUJlhfBeyFdgGmKTo3Al7qR3tBtHCndoQ1hf3pZxQBkLxs1QK
qQy+I8NGChL5Uw1jKkOckKOinlCCyOkJcqGqJks7SSblBwFcIs8H02COCOpjxgO4vqqcuLgiqSr5
oBItptrBn1gxln5ujWTPyBmgnTvqTdyBDFNtOg4wcXOOfSmVAWgsPttG6evg3qcUlJYTaSKxBNzQ
ckOCH1tSGKcMtN/bXcH0+kLgDzC7JD6oMbsd9G9s8FXNajybF9n8UQAlyD0qXYJHsLk30ax3Mtj1
x7t9rnsD+WSkoOKqkbOSorGaBE1dHPDe/+Idt80SvcRwFUOJ0XoCz7SdSlRSimCAycHXw48Y41d4
HqgV13CVnf6uUn6Z2/9qrLznc10eqbzMEuv18ko+Gz1wvEwoQIpw5t3XvmoIDJT1Mb6OHszUi76k
wTIcKA3eQuQ/u2NrrMvuMbSUWfc4fsLQVZJi1kP4K0jsAAF2ucGqr+k3KlZWvnn9APtGc/2aCBYq
EvJjOOUqI548d2E/0+nJM7gJAcR5aykCnHcEp4VV3vVPAN1x7iJNT0Q4/csSiGy4ryIWU9RfHRBy
zSWxgwUk47Ih7GGNkRR/tzVY9zBqAoRX2Zz0XUiaDW1AZYgFXRvHoRoNBqp6OtMH8kDj72TY5A0W
jkRu43aPK1i9QPNmNpdBq3QhLi/0xpwuP0JH8rUvp7zb62vfmU/HZM9IafrBpERczb6OodVWCWgz
zH57xQDQTFlg3vhImharkKRgaBQMASiK+7kD4CysewGTabUYCwGSa0tGDmfTxWw5NFzNiUCdtniq
geRYlFwXJ+Vb3HQDSbnVZkHm4iN5PE10PJ0WgvtJKzjjppDCsatY+8rHuI0eWKCY8d8W2IXPUJnP
h7D4HWPu2hfZjdTrhv95JaLLdPR72yi9ZSavbIHr0+kmfuHGQwwgCUEKpLcfeAqzM6kC7wba81lr
MXyNhlRaiVXh5bFFA0w1peyq4RsiBqOSYIBAcsghPqQqkHt8iIJfous/wQ4dlJDGzBmMisH1VLjA
9abzQMiHuIb26jhtaPQJ1UbEWgd9xAlTMh7tteQ3lx1t0Dblpdlrw/v03FhtsOzNxE/tSlJEATRP
DZoFtRYKQOZsEoPoM1kYniTuhrB5MVENZMpJtG9VuO85OJObcPQveNmhaE95dOxJgRiRUMKbK+tf
xQnQpHbj9BbO2W+GZt1y+UkMfQfi7HZb2BawypRFEIPYut2VXT57ZNDnQIDCSOPjWZI8f+iVdiuj
3hoWgAwx9RbsWO3iGXIB8QsXjdjZVlzVrmMhtm/AhIWvhlgb66VbLkUtvhiP+RAW/31huz/EOeCV
KXjcSuS/zE1FRg7MrREm/T6wZPuYXywQwEOzkA2Qe2JnDGsYHePlffPy7OZ9IxxK6cjTZ2AQ69PY
ktIFiJx2zHr+svspeS99qan0BJU8kJa67rS9AObF9Yae6J3z3C379+2MsmB3B0/Q7K4Muo8ygh2v
U+Xs4XieeuUMamNdfNWFVx0lNH+nUm/+w070gf2zzk7OWhc1w3PK54fStaIJt6TxDXEoiXg+y0bF
2PMW4Xx3J1xGn81EhwjnA5KT+3lmClA9FaJaBVgjulLIToZmRU8hoE5gtHMhI3uv6zKRI4AHZsmw
aN1NUPGUiqvfgmgDt1C4SpmUtOh6j7ZY3F5orS77fktrPLJxN+nJylShRhGiO49PqVojjECODofc
wKtG+WhVl2aRyKmEF51icNRsi4Af+6vWjrKuHmwEkDcmkuuBxX+8qcjyFRPlbYpSPCSEG6XeEO0M
lC1iFHdjdGnQhLUCQzNjQNM8HCYw/Tp0DRB87iwmODhSogqVqeNvWNSxJQ86Xgt4ZHYRmgOgXUj+
2McDjmxdwtHJSTtUwNiSeM9Pdzzgluz92RSOnwzOODbDmB3YrIMpK8Z0Ovar38C3cWByKlmvwpSd
Bg25mX6vJuA8OPnNpQacxhnGhqYUMSzKIBh7/+Pd6dq7giuBaF8KWwwUHmikHUOq9yXwpwkZjbwr
FJYmUJhSa2W/bMuC+UioeZ+aZ55hJM64jBwV209owwqeUIPqFbM6TqdeJN6ufX8KWPCm296YJ6+2
7YlAFnn13wDELDgvroGhbXhZs3/ZUWUt7Aw7rrLfxNnksdsgwYKsQ+ILw5EoTU8XcxC/qQ0Hu12C
qebq2q6f3ur/xIa6p3pE3fGh7pR90u5nlkX0HbY6E6h5yW96GycGxpsfQw0aEVAhvJwQX6S6EVYh
fNuDdbLVDQ7CRv7Y1CaFpXzPU3Grcvh8jo9Mva0JHvnJpGmvO+y86rKsnLl38oRF0jDeJ6ZLUUj4
DjQn+rrvWLyKZgWrjLcIkT1vVH24ZBo3tatW1Y4sD91IUZntaoHisnmHiTzpVAYetvE44ARfa8Cs
T2jmzHPlMidiTJ4HpUi0cm9Wko7I5tI749246rkY/se1fgX3YsXfvDSMaUvKegcqL1ogXIVBP5uo
2KHdhn/6Ux/p6K6cBrU/xx0xNoOfWOlcB/i4vN9Se6QtTNzAHjM67X0IFAtyShZ0xxdlQC23gFVC
T97gyHKXCZfOi2cPrhOglNge+53dyxlXo0eqauLAFUbbmufT7n4kFR5zcj2qvICSd0X9yp7m4zob
pchdRuuwEj0mHZKlLiG+q4UUePO9071RzHaLurM4dYeyaR/o5JhaOzMhvtUgIBp3YvNABEItJrat
ZP/5UE8UPsSPqtYEK/RSm4Lx8J7gi5nqtYDtI72Nod7qimqOo0JG3hk3fEibUlGLyaQCbwFKjEdy
DEsyYn82cAtaRa5O15V/nDM/T+piNZjZIfR38IPQ9Kj3XLywrE0F8ESi2khTRGABDayPuQOpo6mD
qNDE+Bi1hVEnWuksaFdibjAeNbIJ9LIrmzZfh7z8q9x5b3yqafmjCYelUDX93XzPuo/3DjNTmrh/
aL3P/ChFooNnn+YA8JlCKHmy3L3fKJozKrCjQjCLSva4GRImnOL07blPkkYmLvddlwtebKoQxjf0
9hVpJW+mvV5vJeGwYFV6DkNeODRsb/+FDZc9Sq9p6J70vZqBVg7X8yC0l7FhGJCQ85EVAwLCSyqm
fzbahl+HnjyMNNKiisv1pcpGzSylX2AtlETHo6w/N+FplOlI+XeA8znJH5D6fHSKOFbFeX3BOXQj
VkURznonkkn6tqaa7mWbofpNgLeZmNltuDLkxwKVnccvmRVessMFcnVlUk5zASUHC0YHK++dGMr9
eci7wCNyS+ezZIaqOfAnMvl9SUQdxNwnO+y07YdDfwR3/bIZRtAPbeyi3fNSqNVE8oXTY4MtPL3j
K2XZzEmn30e50Wx0RC56LUlofOxfSVO2Y1XnzZRi46Z7aiV/yi1uVMy8wateO4IZ4ORGixozoN9r
lGzsqEAEWV9o4dz3lMSiORsTfjT6IfMs2qSrNcgLO0dcJJ9HHEfCnYiPxV9PFwGYlaleKf/Pl2NZ
hmZvzG89+F8X17L91WPVVjWMBSfz817Hr8NQpJ75sH3L4Gr3itDLFi25af5Gz3Suw0lNUUIyC/NV
viIUJ0p45hyuWiaKwcbgf8q2gdu0Pva+RM1q9TC62u/iXTogLG2QBYJb24ToTtomoLzqIsbWjja6
VQRjY3P6yciIKUtmtYjI29/UstofxsywO9GXS02sHui79STVfHvS+7lEANVYV/3iO2IKOBdrp3aA
RcNWSqJPnv9ahhhAwpvkG5OO52sIAVsE6+lCNrpKliGcs9tRrYh/2YXssi5YqkxEwipsaIS2TtUS
GkescYSvP2hSQTMDzDZF7MDVd1UIUMd5AV8zGzr7zQt+FeyVRT8DSDnIs0nqEVehhwsB3F20PoCm
z+n8NIPVKdxusxfaDX6tGjs4zSPPNCvY5bGpv3LNIvQKcGs2EZrQHrRJREx1moiMzE8R2cfIb/ea
dXStLPS1Ha5CGBRhc00zNK474fsBFRDo2xvS2TGtrCsN7/Am4Q/zll2d+MoHow5aorPAw/c5WCBK
1OHs+1UbuEgEw0SUWCNWgPa+4PcmPteBoLEN05W3OYY13t1ShTF9giiShei69NIssnTcUjb+oojN
TKd3VE8i3KdZ/3/PSplRXUjso9KdA1qgWcuqdCytdnr161104xo0xCW7MB+TPwnVZUrN7PibRdvb
aXRaNZcV9Teu8JSpQek3Di6rHmicBBbhAoJ6A2Z1q1VgwbxqeOu7YjPTnR8qLUi32krODFCaDP6A
Nonr+G/ecTahmaAI4RZbet1hUzBBXFdig47kFhyD1/d2d07SaGkGDRcmHpVN/1OEQA61fBvEQdev
9OiEeuNBl0MT1k3lvuwgYVzYHi368qDSDOKC49FCR1hAeEtxjBAFMTl0xHXUwmU9T5iAsEhTlZ4B
JbvYW37p/MDaOWeytZijTbTLJFHyhXudO2pRuxm5IHqNQpaXW0L3yhLcAZYulrPmGaRCteFbxn06
Hsx8AUjjr2KhrfBEwA7SIbA+yrtn/4byCFWDn0RhxZ0yk2srJ26TDiXvjWH2J9qZX3LMiqD2/1Ga
YbFb8nZHHbYtqIhWjmRqWia+O7Sw2mA+7BNcByCvkF1vbt39X+oa411bkSTp94jrUbn0xyqHIlvM
A6EoqT0Dx0H/LqJuicdW+TSdVAAbBHHZZKuG5tgC+YTE8xvUDfD4YFCutIqZL8MfNTOhaMni+Uhp
7th5WPun8grYopTnps25gQzbmuiBO+0j2ex4rqkbTf1aKJTEOjr43Rfq7s88LGoKtmU4xG1b0idH
GpRvnOCK3rSoafSxFhAdlMIQd6WzXdjSPNYhgrvicn/ySVtRMrKUlvTGYMjjGdKhEtku3D71xV+i
DM/tAl2sGS0BUKksYs99qxiuK5crj3ZAckRH50J9puVtIdFR1goq0cNBl4wpZg97Hg/8yjBhXFWz
qAztebWlSDSzh+82OXkvhq1lUWlbpvWBU//+LGJynnfuHUFxCyU2SI5Ms3JuQQZgZ/LonMMbCvwa
1uqq6RPaWMJLzyrUPcYD915deNDiZaqOJv2KEbk2WvvLlKDy32yiDJszrbMbCcR1vCnEs89iTqHV
jWxmVxxuwbwsWb6h2Ff7ifrnq4MJ4YEBJiH0xH/DCXUa+TDMiUfmtFd8cz7g42VCGy3ffTgBx3sM
/pJn5MDvyciU68Wjkke4DTDR/coR6g4FHdRqHE6doBrsOLYce7jfqiWCY8m2XU6AKL3VNUDmTsCE
GvBnBTkTfSJNvMJpRIga0EhbhI6uNTTHU5CvnBrHcBQSMej1u1uwPAR4QDboTu2JpME5BDk+K4Rb
S36+mDyL5eBZqCTGzcMgDv240Zjyhx3edKY8uqJ9abVo13g4JUi6oof13gCuycm1huJ9WX1Ac+p2
PhLcSmDMplJzAZMjQR5l1YAKPUdtqWKdggc05CzWJuWKgPlI9GuKRvO7ilsmd7IDk5oCH7HdS9kT
wjEIC0mKK6JAUI1zhmpalKnYqwW40UTHzRxxIXFv1UZW+FwlB8Nda6K50LxvQQsl+DUEMThtApYq
1LYcAnFAwBBa4hSWUTxPGJw3nfq08QQj6rSV5uJYDGu5iHyNWE2LN1DBe7QKghROo98kb37Ud3GY
PKn/I7lh3+4AgHm6CwbW1D44bFDAgMcNcoisMLHw/Hf9nNUM5pW3bZlK3FuXLTnInzqf/Pt3R9Tc
tp4rhrWvG5wqJ0xbeEFaHKB4Rmc0G5tZ4N8zveZHLZ0CG71SQGkDLWtCstuZt1iz4OXYPCGlpEyH
4f5A6vZosvLoef52zvLCyTGDEvvyzDCvtS7jYPDzmf5J1aP1O3tCYn3EoLNHq6iZMaQEAzT+iDvM
F5naAL1fGr1avwpUWwrUDpWPOkNPRzyY3L2udbAgB2dA5o1hOXTw+fhmoahU5E3gPVIiF8P6zGbv
0wb8iMtDHckTA7CCIWm4gGgJ2s+8Wj7YAoS+dBAUqNweZtLbpNRmczYwnJeLllzyCAAAWEM3F6CI
bIWf1Imgndd+a+OfcigicG+nHnkVDL0FsRpXkY+vy0qE6yV3uka5i6iGEH12zRsayko7PKeJnaKs
Bm25rfjedquv8eqonXz2q2ohK8hlmoeZPdKjTi4rHMtiYYvHQJuuN7qU6xm1EAbsu+WjC0JILtBZ
6tz2XaIk2LS6TOunnuyeXNUVqheqkvPVg3Le0w/WySvEfNnS5nXYpz5JNLADk8XR86UodU+irm+m
7/uY81LaGr1EKibm/lYd7GHnNGvOG6hsR5jqYkORKF8Kxmz39XmjXdcp0qI2PrgGlyGO3y/810nP
EG9py+IuGO0VrL6XI7tcpaB15TPaqzuHtCeyv8tzffVCSM1XklqRkaFd1zJQarJcTeSQ26Gl79M9
aDnM27Dvh7XO/WeT4K9iNrMG3pYJgRa0yOIZ0HaIL6yLnrtMks4wPgbRsXAgLvbNsI2iOVnRqcYw
8qYm3QKjuMv5u5AF8n6G1H+4fIsz3QZ6GPicMB98L1Urpeg/8bfJIa3u2p6PrW+nkZRKR/dmCoum
vSVS0e6EELYYQMHi0sZxN5fKdkh5lkkFXPP2kaEWlwVknmVpxBc6Air1XkSlQ5jWkZXFvrhlADH5
fJhx9RHh6Ha5R8PO2x4YwFxiO7S9KsbzKkCrRRVu8q/9nd1IVQ1dUknivumv0ykkYbxT+zxHmmGa
cSmJUMwTgMSdCUGh6JETL4ca1sJx9KDLLC4YMxf3w1s5S40cJQsJCKpKCyaNLubsn02jTWXUEdjo
t7Su0gRjqArTKQsAbgconTzCBaJOKo74XV1ljVz2+BGs3yJaIuTm5dPh/q1xNGlhFQlNmJTBKkaG
9bSiTzt8Ptmd6QaHfKSYD3WDh3VLsF6aZ3i3rax+TIpc4FNStZt2SjzJ9rUYo224wm9KOEDy9tZf
0lYBPIO2PEAgwr5X6uZzRsYI9O7tLW5cq3fd9XXEU6adr9QOkKTI9gG/ice6Db5rYmRhVPDtle6j
6KmpE3bo84kNrzQgqUxK3Y8DrI0ghpHMUzYZB+wUJ0hHpC3XYxMWIfJZub1kT2d0v4x+lgl/nK0J
7TBHDYHI8oqIkyZzni8w9uLy/DyUmrrYJxrDEz290TPhAILUAol04JUMH9WQsE7DQvUp4nehDkAW
ktNfm1P/7PRKlsLoSo18h+jSGTh2XFrMgGiDNqDNUMIXt5aW2oYSIXbhdwo3F+tR+CZERWbX7xB3
+Oyaa7zWBYxfwM8/wN78n38gqhkS5UuD61VlSM3o8DhEyyRjG+4BbtOHnJKq5tD/f9Xird7fK+Tv
7i6zdyIrXLNJ7WKR2YXxilt9BMX1LVHgAqqeba0dP8FNBzJVKqsDp/vP+8j0m9fxu/Bkyd+em/Xv
hOKTidBRM6lRxzu28tktnbTqHEDpM/i+pw/JAX+legTq52OdqRHja9MAHNA5QEN3WpN0Hj9ohEjY
b1bRbIi5AwuruO8aHLA2lw5JUZ6Yi2EuBDEiwJ+xbBa8/yAE6Y0dWN2BPbtXvNSYINBlrG+EvuJ/
5eLGxhBij0N2Nif/icjKiSTn8X8ruzbO4sGVmkkeGOgtFpL41WzSP/6a42qFgpsLU0wdEMBIWIUR
z7QBYMW/2vGSKVQ7MmRnm425H5beui/pzA3wUCeqHdQEpw15f/PDXctD5+Ply8kaVRMrSIgCz9M5
X2y6Fch58q7X/zzroHrNvqgHW0wgp0m0NptJAyjt973OHRC751Jf+9L1jbwj15jijHKh3E+6F+vI
iILoX2SWgSS+bImvLa1gPtcHk5skR88JedYNT9Nb5TowApeBlRtUeluWYvjJ3hQjeZ60podYm8p2
3BQ9X6J50nh1cgBHkcQSuuxQxm44lEHMMSbnHM319iV0O5gQXfaEekHV6qEH7Rvoi7kv4bevrpkp
RbAtnc0v2qQJ+Oisl53hkeHP5Eft7vOwxMoYcF9b089jQfq9taScsBOCEgrN4Q0mRSqUnpH3Rhd9
nrSnftEi6W56xplH97X+KHcpnyB4Cl/wcoVi5uG2kB3Q6EhtGTy6sPa20XUdStSLqKtEmoYeBmXC
Vxz+qDuP0uDtO1xLEvazDOemXa4MMhmYcSXc0OZ0ul8gg75sHG5mKNgJQsUnhHn3F45l5BEidhjk
pmJCFeFpLaes3tYP5BJWWCxb2LaGTLlV+jgL5ACgqvWpEw/S5VhMrzseCysWMg13QG3k3l34ugzd
7kRz60E07udgZfcwKmYoU2hcnef8LOm+QfQEjnbAWkHLUE4OUoIzNdsdDCY/91tjwz3ItU2xRSCt
jP38XfQ8MU989sl2txM6DSQFZLcF4RGtvXXnx8Z4Pfz9U9KhW8gLv0CBeSi4jYtlNMj4s49vBm5U
vVRuDB9h4l3wRpKgxEMESmzAbb+vlMBYgbonWay2Q+hZexPZY0YH80jeJ2g8fhIVHkMcADF+DKB4
CaMQeh8EbOR36Xt/mhgKF/vCyTfMAWvtgI4dFdo/lzjPXu6ixfpfA3BywGyfnRqp5Kv0Nq7oxiuj
e+1ZVJEAyfD2+Uz+2C4LDyMbesKMvhAxKINiqRaWmIKvLDMXAn95dvTaskGMkrtBkYaJjqq5g7na
KXG3siAeoZNsVKoys4JcADJvaUvO2H7kMEIZSy0AHyKpUjU1FIRvFmdA58j9rKUOuC8lprzVeFhe
/zY5Aw3GVMCKzxFvkf0QBy1Fh2ZoLvMGeL605H1KIRPCcFx2FBusO48jLB6+mnoCiLhqRtdQyDy3
hLnhQxrryt4DU9BupuOkvPd/UO6+MzdRf+GBrE9jemkyUaV2IpWSySApeVVz5WQ7S1SquZjAqOAB
CaqSq1KafUbXCWW7D/2wKpj00I4Z/BOS1QlXMeC1sbQ5WC+32WPr6gcslfwvOg7ZSLWk4GzbcXXo
9BCUWjtNSOwvIYiD16kq/OEyz6Sagh21p7tctx/O3jG+5hZDui3S0mtldOjTq/2gRANTk2yYsabz
w5GZZEyNcTMejdj1hASugF7MUmwOmut4xPYyYTvmnjShnN6FSz+hDu+lY47932+br+rHi4bEMahb
kA+z7YOxAKVRGLcVcoA+zuSaij8gDq/4esox0bQDgady/1yZsVqp8XU/IpulrpYiBB0nXrDK6wFJ
iMfwYIXbEwUxYhV6ANJKOrhkrur66Jn3ebjA4z+anpynbd5fOMJHe1QsdFMkBPgkHr7udN5mZVk5
5vQ9qM4vUdRe0TErNZsoy66lGVT0yblXeYlVMY7E4TEFgSzagNleCmNbdQ+FrQ/DdmVQrGVLBDGk
azb1i8ybpM0UPdJw/6St0McKBc2ra0FIjI2wbbCWLeFFWmFRjoZmioyItD8WjptOLHSgC7yaCULv
CawD0d02Re+oJn3fnTCERU+fw+MuFb4h9Ii1y+aC2Fh31ewATyDx+g4pO0gSR4jtAXyxm/drQKaR
O+iN2A8lOw6i6opDW1aU/7GrTYjr4Ku9TYnhwUwRfA+tf8Nh9/jsHdMOH7BRvNursL7A4VOS5uvp
l6FgGmn2WOPFMBQo54Od3TiQKQpLc0upFdwszkmp4Ng0S08ysB+QI/z48tt06Ru8/94veKSA0qs8
rs0my8ZljnDQc9bLVHFQHGpg32h/Xyt2X23tBYGK9QMB+uEe7t9Uc98DkjBjNN6bTYtn377A6pDK
vvqlKdDpB86DN/sowdVbO6qbGUPHKCHmsBpeF0m6TgfBEUGj40wLV65+H5w/VF48iyJ6L4Oy0TVA
mcQztjwQLWeaQrQun6v/qN4vX4YSbZn5Kym3/6Zv75fn46gZoA70oNjuTJuagstlLvgoBDFEaJkU
4aiL793dngvNlqdL9d/e6pgDRpQNxawnEeEFxtrQfXJl6z1xp+vXdLqX9nlLX+/2cmY+06o6tra7
CCNg1tPldA0i4CGZ2YnjmD1LSfHz5X+Cpo5WmGySe1Si8JjrdzsHsxUSo9bMzPf1vyPDBcjWaIVD
BK8GYb+Jpvo59WsZLOn85SsVTCXkNao9ZcilZYOSRiQQJqibepKXANLpMxN7iCn3GQKjnnvV9VvM
CnXkw/dr+7ohmnc02fJwSUH34fc5mNHhnxpL07ZgccCjFOt47aww97V+Kadl3fQFZGicJ8hbG24L
B+Oxy1Jmkh5ft8ap6tPX1Gp8BBJGVNvD0uVWt3RANR3KbfFlmcrExq00kZP4lhpjue91vnIBA2Rw
2mj+75PqNejj3oTGaKBwx95/wS0NaIIMkRZEqID3PRAcJlDoJO6+Z1138iFfF+XgOlnHbNEsMnDl
0/Pp09+ntoib5tH5xuKueFXe4a8Bd35JanoXiePFT9ZGiFs351Fo3pvenvgluwdf6aQFhaEDIYM1
Qd+LvrMkG4/tycMEpLYdOSYY/ORWhcz29i7aPUjFvKdCgymomZ6IYDO16ZB1CFAcirHNmrTYqkN5
K4xxXmKPn+A/J2phoz0/wyg/IO2cA7jIOzHt2Spa5VlJXmQdadk8S6/uNocbJy0VQFXoaoeUxi3G
kDkfoZQL/6L4zaALP324/U3ZySMcfFzNOAQ17vBwz+TczMdbfHZObBmWOHDnPNGcBvyfX+wc9bH+
pk/WP06grSpcamy51f5YZRezNX6yIBdVxEIxLtUgRwtSK+3VPT4oZyHiMrNon1agnodWXFn2WR7R
VUdq1MZ1pzrN8kxytKrG9OR0pPaSYf+y1PTE5oN2teMZaPOkwTXuo9s9UdP4i4BU96+GA/tYK9xO
p/aJLnCBAWRXmLS7R2IAFTpo2cMD2HH+2x5BcAhekpZ+tLvmBQQISoqAjg9XdglFT7REBKh+0CZy
cys0cZ+S7A2ig2sfyTTnnsq022Cvj5yRip0OJtb2Qb1mtVNXaSchXF5zlOtpviMRNIdpds1TaIZh
ocGHt7vAEO3hvjOfRzbMMpf0/Ce/kEq2zGYc6ke6EUUN1c1GfNiG+axznBFuk1YkTpr8Y0xDxq7z
v6lPvre5mEx5qFREX67xNP5nd0bLISv3M80EMceXGNLRVl7VHbiOQievFd3ZZazomqkipqMFj/wd
Gtcdl5icIaiPwFKqQLEsIfln6p1wtYCrMMQaqpyBnJJjmo9EL0+ChYXXtzgMR5syMXkOk1hiZhHE
sA78FGUASDy/WTJOsQsriYqSRocHIHf7lVjXjwgpHV0z+6CuSEcazoXLVU83KQhuCDUZ6+5IeORp
iCiv6z94CPCfLKznlv1QOsHkENmOocDPq7GTegdYvUUSgEwQZEgd9g9diP6WajSUYiktNuVLngMC
Gh45+Lh+usbxJRZPfqzq/pd5o2uxdAzHPS16NoFq5TAxlmzwYmAIAAewj+miNuvzeIgiP6vF0SfG
DtoUm6L6boQWtBbQ/0kUmhPh3KEzPQdKP6q/V27HgrulA7bL9SIfd4lxJBPxmr4UvfP0NufXuaHX
nnJoqEu492moUXNPv7cN2QF17G7Fw7/7buET/wBV+mtUVd9P2Zd/SmA3IOvqOXBNIwv2ZWLoemIG
UoU7OcZ/GsDOcmYNiiPueQqh/WcDYpNU4F0YXkgahBeufTHPjrAqEyWsYbTWytN5jPXr3aNPkH04
/pOHH18A7rSHaZkQJQxYrzdSODyORqwrnUGJxOILgXNTlJsEpcDfUWcq1WMM61b80asUh5AYcY8a
VTcItt0Le/Mz6f2JILIIpT7SiJ2gx/ODvA0YZ2MDesCXoz4yKWSUguIZiMGZWZr3wJWyImGRyJ8y
Y9JZOJ54DfGxYIohb+WQzzI5Qo/8qY5LATAaP7VC/mjmJ8Hjv3/oD7vACRP/rJ0vJYCoKW5asidb
8mnGBTuu6F+YCAHInG8yiklcwypeG62orgfkJb4qr1dbQaf0szl4DVwAiCB+Qf0LqBd2zdRAlejo
YLfK3Sx3NiqKhTh6fhvBjb09grCvgVnNxnrqL2KgkqGEEny3kUK/1NgQLv3GNwxI2zcELkkziO7w
GKR8nG7buXuKOrXd++qO5j9r58ITLyewJdmgL6+w7eZGFILksY/RR6zv4xngOv/esqjPBfucjLlr
hVVPqID1KleyIbkiwIwY8TNwjnA8C1/d9/r3rgmMbmO5ukdXg5gD/rTTKm6BIKTC/YupE5HM63EN
pFbNvHjBr+s0YFvnntAHrZ0bKVYaIMSS4iWl9wQPcegTo6z/MHO7s+GTxGOOnIZgf1aG/+gmOncO
/hHlFrpMBEK2Ba4AF4Ys/ONV4pg9US4VwvRCmzyGzcfOXi/SvYQdJT8mAFcvdaAH2xQ0zh/ETb4V
SxklvcL2x8c2L7qB97CVmxRm4srQt6ZlILefU1X/DvnTQ3CxEfAVwugheHme41Nm03aC0W4A0ESa
kbovSI2deCJxpGerBAKztdKNVjwvN3h4blTs3eIkaVwH1yh0pcNKNFqpiyfFSStGLufapIBNLgWD
q3ARJGseTHnXPGZyR0qJpmL+VF9ji8ZXpHm30m3V1UtDk9E0ydR1WPtmsoG5a0jhXEha8YyCFWqg
z4tJ7W0+9fIRuW2xlE4ZWQ7pAMr8zw/4+XDYemGGWwce0igSpZfB1gzmJVXWFPeBP/yKVZMyny3G
T/9D5m7umaFSOnbmGDVUaeS2IAXuv54paOvrs5NU0A3BbXGkmrss5k5RosP11CP4iJbY5DXpLr+R
7XoUp6z6aUitHlPW/juR+rE0J3li23giSbzY56dfTjNCUJaqb4NcOfL0nxYFA4jJUIf1iC7+xZIk
sSfor5oBe+1gpNWkWWxapxf2qLkcWYGX5zCaEhhT5to55UvRiudXfQbYcKqS41PmhJCF2yJKAX0u
BO9P34IufNmvV03237VsrWN7/2hv//P1BkIvXcW9ye5pvss8D8msKobzGEKAYDL/qc6yqlNzLhSu
XnmTyFEb3Hr+Gl/BkgI6Rzz3m0wFKSnIKLXxA+KsQ6qn0Bp7zg5to3Mbodci6gHjZjPfIzhNjmgA
BJ54uVQAXfndsLR57qW0Wm1KQiBBot9+bor3PbcXTXwo6XOzJLBrE2EodspzH1pMs6nBTK7Hv5MH
NluOKwZuGA5n1CfQo5jdGtQzZNFce7gNVO/2/7hc+cfrj1Ul2WR/zcpxzOEGNbUf0mnlJhNfREha
Hytwj1Q+qvj1kYmj4pOLpdRmZ+vbEU1MUGeX0ceXttchbZfj8WETOqg37zxXnKD3T5i5gqpwNWgN
n0fRrXkaQJgxGelMcryFJZT+xhxAf8hXP1oCg5c/BcGp++xaaRxEYWlEUgtzrO7FPSIIoc8R9HKB
DGQAuSeIMsrgu+lK8piaTIih5HdoKxlqGiS98dItzI6ZAkxMBSJPjubUyRzRKbHKY23C6hvZaxms
zVA0XO+mBad6sQNJKiRwhFhvJ0iq596FMeR9TOAqqbE70ZwWqp82aOycmnkanMYIMJykgzz9mFnB
laH9a+4VMtFsaFhD12Te4aoPU7HdsmJE4D6Anfui3kEZQHPTswwWVZx4GFvU+xSiWjI3HhMBg1e7
C2tHm7Jsov71L0rDLmffhCRm01xdJoMpy/x99vw7Nw2Hk+eKjoMvszhllGE9qRlzrX/KHZXBP4Tq
cMDvANHjpvAXvILy7cLWEOVhn6lW67I6y4jhmWSgXGFss/njBkrkbjzLQB85EFXdr26RwgbB0kd5
pCEQc7xzZm9LK0ulY1G4CBM5elS92VpBZPWE9cpSeidFzxh2Yg0/Lz1aYuOgCBKGsPdjK471cAgf
kdr5ASpIoBMNHmaoRw5BcW2NkDXc22VuLE5ANCgP70nSKMHZ5nWeSM1YRP9mnnqHerkUo4MDLGEa
gbY5bWW+sTHBeYtXHcumU//oIlnJc5HvYjJ5SuRLoMfJhabEsdWK75jJmkPhSmg7GTgaYj4ginPa
e/SX3UeKxKuwuD/7SL6hGWk5FfAXkyvxPh3kEMH3BefM9EseLG6gUAihELLFzu8kEz9Lghb3zJYg
PwygOqF/AGQHi/zHYIVlpABTOkMxGetQYrPxLPl2p1QY7IIR3fyfYtS6ZcEU+BNshU+QB5gN1Vb7
PNRH4W91izBFwcG5Kj6AYqNfWfYQDTFb/62+eLKtNOdMUb9uwFr8K3NKXwBvPxQN6xg4qIE/pCCf
PUqA4wlo0E1zkFLVyqX0xCMLSsnNvQjumhGpZi9J2qjd1ww0dnaWL3OzlNYtx7TW371eeUUeNIhj
pyChXtYXiAIJFp6Kuk50W+dx7t9dFPPQAWoi/3RdCRYWWOmOTachV4noDdxb2zKKrzYkjyaXfMCJ
nyHz5jxeCX2FKFvO6nQgUHDe5ohDaIoMHW0dS6/DWwRvKrjOFj+dsMCvqHicW2dZ4SToF4N/oNv1
ejjU0JNLGe4KjlqcfEwmA8EcAs8VRg4jBpjlV0OPHZt55DlfZPcaOdWoX1t2Kh0enUHHsIWgrimC
TNPEB6/TW0VoNQxo3qVTYhdrEJxXPSEjmfE0GqJc/ciMIN7VJ9nBR7p/rbpWO3H0iyn+KYuORkYo
3LqVwV3Pn9rAMVvAd5URiek2O5w2IcAlj+ghZ/k+LsfCXLa6RTcDmgOX3L0tilr6o7Mmcp99CRG/
vabgYVsVLJfu9T7lcC685TBG0nKw7a7ITbBJvmgWWFrybBCZDaNd57gDf9kzUAh1CL59u1pu4/Vc
QmRUdg3GsuDj41j10amnNnLEuNdPow7Y21Ab0h2uyN3SoDMT4/NJWeSBI6+IM448dwkLkluohify
AL88If8Px8x3Ho2KUaWNkTLrUbvJRPYr0b3CdHszJq5Z6oRdSjUKmnHVvqtx8ixR/r6A3gvKAHRR
SjuzCPdSx/NAOPRH/NJuqruqa61GbiM/vpTnuFpwdiNk52/dKS4JiRVHCD2KLI4w85QHSZ8E0mn3
g/676NFbdTxA2tAbKk+kLpup3+QS371CAMmh6qAvAn4qw6KqHZiFwJN7PlQ1mIm3M8BoYFvpQWdH
aaT5ixn8GEJ65zREpyKi/T4CV/nk0ipF8Nb6Dp4+284hChbM/VpzLloVia2LAwZ4u9ISjy511Tfr
XbdT8ovkks405g8y29bFHrlh776PSeYomKOnPXUkkHMgMwz0Lro9AgNPkL6iF7sGUYqpwvLp2aJw
ZQ+E6dwHE8pmJ1CL7Aa/3DA7FOFVLFXv5SLyqWj9kysUNKAB1BRDUgIKpf5AVuNqR+XnjfBJwukL
/H5WJ5MH2E10bQAjapDbhiboIeb2w0CbuuH4Tmxe71QKOYQMTvfg4zN/w9dhct5qU8MkBnjNkJ/K
pHlhhojDHQugXUhnEctsN09oezACXgFXw45Si6GPPFISHxxr0QgwJ6euSkfsssggTEiLgmPqqKq/
eNvBbhevZzrTwsiYOb3kZ3Ysd3NRVKbCQv8jNC42N4j3uV3chLj7mpoKEPV/mDxaKdQl9JeRJ9HK
d1/OQdDBJYWO4iJwEz93xTgzUUSwh9fJ5UWXPiyi0KG7FGt9KkXq0P3GHfD59E0guPC7NWyOcgtP
hZmmL5AMg0aWUNhXfbB89u7tXgfePQOFzEk98lKEG5wFmvZXc8qLrkubyLFBYbfgmdHkBAfLndjr
e7bAle3WByDFXA9HJnvX/jROx9G0lTltWTYTvh1ncwTZRN3NggoLXBBMCXfUdKIs/iFJbIwMuR9l
bFDlevPx9qrNPXDAPg4/xoTv/n65tuykiS266vK2AjD+XQB9boOSvyEMkAG8KfQ9HE5ZuZ9exzfS
a842AS6n184+mFtKdQcA6yBsrNPq/3cju7NagGSb67y3H8r5Qti6VX7EqZucqsmLkxo1IGjRvjyM
bvBuGWcvG5GFJUoQJ2OEmlLzJJOXM2KJ15A8ElGZZaUc6SqsoKsCLPN/D0JhFS123lBSDV8y+KJH
bYaZtgkiEKWNR1Mo/de6gb8NqiYeerHQ1+MtZZBcSL3ZQQnv6fUHp+b9+Sr1g0D+fBKRzkvu4yM0
/NRgX+GYSaMZ4rTPZ11vdSuorjopuWyxamLiel8/fVuapz82HubKmGbpQTBNL8lptsBxetvz4VSI
4AdrobCbKtuoug7yGyhxUsVRwRU9jGM75O7gERmJdZOxGNK1yT8cZy81cVvPGWW96lFUHXun98bo
ogjRZQ2pETO+x5vysCsqG7DCRog2AuwauvbJnISvWWNk8EfH7HWlP4xjmErahAkoX+hLaSsQSbtc
sLttcS138VVnhIc6BgAxr5ft4IMFm4BKnUUcaFIr4+SR/4p5+hZJa3KwQmlLbl+5jMM0mepag5U1
7jw4OcNDXOEttUHQTFGmrNiHgceTk4IjKvTGgcMM1iGTi4S18lO9QTsySkjSvNca2W138yWPSkCV
/7pxcFuDViCWgau5yAdBJcFfVk3W7zsZAH3rxEXvaA+hlxWM6BoxAfR367TvavJBeibolv7DERr2
2/MROYnpFDY7grYxQJ6XALjKDrWFrQnVIW5xjRqepNA6jqOSh6FmDsYNanh6dN6gA38sm27FyNi5
6Z76Ek0i7hPfKs47cvcku2VkiY6Yg54zlclaTvXDrWArgCmJRb0+y1e/HPq+2qHrhuJb3ghteQqv
qoJduGCkDBljF3tbAPjQrKIkV2N9JUdDAM/+9t/M8k7sxQid1fSb4GGFgexbdsUqpnkxCLIZTDbG
Mit7o4ejnWgoPyLYJ5wggcVoQJvNKLkXkMGpWD/WJn4ffCbNJChqb4z/yKc3xcecXyHi3vOxO+V1
CdpOfomuDspyDEMgET7o17TaB398qy1l1xsCDCJBWwCoBg+r/JK6dxdRspXMQbghjiNH96bKAXP8
PijS9tagROJkTNgF7XY59Yt4tPtmbtSlhWXy2aFZcSneUgG0r5reA7Sbvi61vJsAD2I+QrY9rQD+
huOs4ffGTbHKuNwMyFoEWmeZXis0AGkYAYc3btVBmy3wc82DOixO/ILdxr3doN0JrtHRhy8a9702
bbAztH1KphvjK47uTb7J4m2M7TopVnCu/h8OlzA7NNxhg+rAKjTZ7KnII8pOeY2NT1JinN8K9Qhf
cL8IgiqKEXrvSpe3D9eywWk/jyHPnBx3AeJ04/X7qltgpR3cb+P2Y+M9H/izhm4Xwkep7LfGnzxR
LhoduvnAafKKVSvRFmld2gw1a+oqJwfVnuJjqtOalNxqavYX1kF9fqw222a0FHq2GhJMncncMOmN
eEh9yqa5x+WwtpP78THI9tY2TRk2TLSPQTMKtaOMrCfPnPsa03kv5imD0bnl0eXJ7XhkZT4fDqNy
L+UZ4YVIpeX5ulzksZlbHqdttbeG9nCPOfpM8FMH3kvNMLaR8M1toCOvkrxAusDPSkTtWLs4Uuqn
0hOQfZ1ua5LPRzqyf7n+ZvqfQYIJS1ekjetrBNtYGjIU3XoN0201l6dqkJ+5UeX4/2HHqjvCtXCw
dR+csjy/YZsKGobBVaoj/mjAGL1hb2iQNRnuuGvyQWSWDroVd6A2lo8U9tDpev0Nt4zC0JqRD1Dh
CvUble16gmXyP8w7cDDXzULKnHSJwWXMvF3Ndb3/nSM/xSeoo5Na5he2IHB/Ovj2T3j1FPSSEJbd
H1+6w4ijvoNWWKp14xTlPk6+fuS2gH8rx2IY1n/2aw9v6qC99HE8bd0JYpsm6ln+qm5Bg21oXdzw
sCr6wEGnle4xpxZfDXgw6SesjLFuNnxoct5Hv3QcHo2x5QMCcMHN23MlwSxOirizjYKUayOxMHMq
BiBCFl2ajsPLm2GJOJlrglc3Tdar3u8PG6MEGAtJfb2J/6HAPEw/xeNIpaNz4bGy7pBhIp9evSYk
UeNhKFhr7OmXffsxJeKel9j19zDCXUGnrtOcNcfojuKQFRWaY6hDkSDVnG1JvhFpdLHJKEjB+lC0
EV/lT0EBzrtXSzHzrMya1yLsKeKFPvaKeFZlBZZxTwKzklsdJI/SZHS4tcueDalESX6xh7l2rQ1O
7TCZm/IrmM81Jyj7NCb5n9deBcbhPfsWNU6Zg92N3mU3U2qavkuRTyVPW7iGB4DpejMaG76i04B/
BPjW0Tddl7aUAyotkUmXy13E6FkHv8/hr6M0jSeVExG1gwkMII76hx7DIlohQzWnAfnWpa/5EJc1
lAHr1ZSD6QA07Y7JZjGyg+LOUlDSvXIIsHT5uxl3rUKgvSUKe6ifOFgstLLinToBHcQYXgW895/E
2dHFCq/Kst1IBsBAlrEXTPGO3LksTg3cIrYWLkbGM28N6XqHuHm86Jc/z/zfDyNPUkOEGFTFiop5
vPVbX+mYzWk4RZsqL7A6fJMmOsdaGh6Y+jTe4vLbfgqs2en8b5v2pkdl/+5uu82IUcvz+4DoeOoB
Bm63toeQNFJiHNDUgUNoUKJmDWmNh3T6jSvlCYNu8KrNGbwvrW3iy9OYv7etwGx3x5SibtZCmOai
FgEPN5+ehELXl1XwpanazGBHWSBOtae9cbv0dVCbXxkHXNyqBcZlm6X+B+7zI3jpoo9Za1UEQIQQ
Jv3cCZwNaGh/bl35qt/5v7sWRP2iRQ+t55jpxOj8zepWSVWO2XkbD6gj1uxNC45c0eAVh057idXq
aTd9zzJ81r8rRYonXSPyRGHhNBIBIBoqWnl4SZK88M5fDaQ0SPn5dm4bCwfjdni2UIjFOl4Tpr7w
MbKKte5oNRDhpa82nBkQOxt783mroKRlEB4/v1eImQEG4Go80AlMRhxsK2WafFfcF1U7BgDtyVsT
6Pw5ClNpVH2xPIYn/qhKkif4RhDTPTQqzBs/jP+PAKcXNPaEOOf0CINFL9NkNdlZDR1mOgz61HfW
AjoV2oBI3q/tsYihcNyInDbxn8rP44WNb4rxn2nqI6nNKEUDk8SI9rj+dLNyyjLGmo0S3LKvn+5c
y5kiZiPU8rwrSd+qjTmdboEZtVMqAmFZQx68Krii+WUyGDz2qR1w0sjTBPW3KS6BTsbBZmKR5/vN
L7xb0oAo7g2mNEDYZjWSPGqutTdRH9Rsc308Y6b2UdP0RoEbnFkcDeotZIl89c8uhhzqFVZB6+21
oBdogNFIZqSieZhbdKarXqxtxG57h2qoqOeF07yhFeVB1oapcTsCb72MTRiWvw0Ufitthwx2hC4b
ZFP7H73W7MVzb+CVBeIGOlDwUVUSPkhfFjogsMFyu0gHZEGJOZxy3wpt0MS6GYusx+JBLQPcBj3X
dYrwWWo2Aow75c0NmhQg/eDIO0uFDozOun0Qvk3ByhA9UcdN2qvgojT2cJjXzbz0z4TBZJpQvG+N
UYf43JdGcEp55XifrcaiXzxtzybmOsrEWjT83dIgnWSHfEIHi/vvepuJaWitf1E5yA4BXTgKFt3X
sv9Zjwq6S7o7hU7m+DQcWxFoRQhbSivFXFbF/HqGZ8yls6HCQryP0pF+bzBc3l6tnSC7w0Cjn2Gt
pu97193PHfX7sOlJKncSPaN24bf9CeKcT1/MXUQfogFfcrt5Y2M4Oqw1KOzqwGFz5aQ1gynqrhMy
GGwGFGMQXEKSUTvZEOTHb+u3QrKYtaSFYKgsLWwAL4riw8JGRP/cYqBfen9TkFRgJb7LpsY08GUV
PRcvaI1DeZVCNz68jbdVOtlxMLMV+sU9/qhAEaaEyfBMMBac3f0vqZAHmJPDLKGEGp1DNry8TQTD
sDoQ1cmDn63wS/7M31dJRy4C1/AHurPzpj3DZR8o1o9wuzdOY+TrmEEbWnIwWa4XZpre+eHJGvPN
gcHiIw5XNGU71tlgHbpaCmXCD+Z0cL33MJX9PdVNAim/eFZ5n3xfOTV9s/FN2Z00MXWUXfoa37UW
NnDrHcGyzp3GOQml4lXAEJ2eqwjieN95DKdg8qqiVIPVdVRfWM+BDNNysjACz+vkEPIBqOWhR4yL
mjYdTqHcjSd1QVEBOafzcnonGpNs6+tqN9CeMd+4TAMto2GkWhYPigEcEZigBjWJgPYICyCJ4pTC
QeuSkVuETEFTk1Bq+bJpoX9O4ceXF4XNIY7WYYBKBWluA0wJ/H6NI3xuOJwYl1poMZSxsSsIAlgV
rR82B000yA7qLb/JdDDpvQ++K8xiY0tcYyWy9A+Y5NPvnsTkrVryM6oF2/q82/51O6WhDTQ5w9df
yXw5MNpRZAhpI398uctVYZhZpQErtILE0FuzdjpWepFShw70a7kENXpY1Vo7W0FRjoRCJrCQQZBg
pgr+yJjvkcWWGGDtE/5TaNwI7Ui5JdaU/evRahxQP2JlKsSGKvkUL5P7Dis4D/MmR1xAGvc27bVR
53a/0RVgsKANiEEqcEPD16UPMDBw7KXerdNi4m3dJdhfiTMb9+ooY+0RRWu/Wfy2BO0R67humQOR
ddC5AB/QeO6nGRUcXiZ6ENeDkW/rFat5lCfiegQIjY/5NT2QKHZs7hdJFHTG967DP3J7jk+vzzI9
NqApDiZ3Q170uU2I8dascmcaj0rLy3qxXQ4gnASNsPE2eI+BwVhyRwOCf4ZoTx3X56IjliWJo4l2
MtBpEWL2KWv+eo00lIIuxp0V/zwzNPZpC971t8KnZ9RaTVYjkK9Wdrpr0ldx4z3Nfrs2aIoyS8fY
PXq5ltVmoxidL37n9USxxscdeVGHIwOEA2S/PiaQWevVaYoYiD4GP/WyAyofQBS1EhR7WsqAaw2Z
0sdqfMMsK6hRnzysuqd1Kqe/jzy7GHY2fipLxxDIDFbWoSN4aMnXLamBvzRkep5II5CEHYOiAnsQ
C86ld1nswB0P2Qd5HzTkpob6nFalpC/LTBT4yyidrwEaILhkFdxJ2RbUrlAFgWDH6h3Hq1C8LxdI
TLIAhLY1eZQgggkIj6iAF5uKUUICPAPfRvJFuzUWLKHJFnBLQoehwe0ezo+pK2FGJZFyyqEh9KtJ
M5xISehAXYCwEBZH0EtL2C0ZFPG5NKudHDFKR0FdMsxvk4/DwT6YWcgwfsW025ShlsIQruNMwCUH
H2q/L+e0QXNVHZQZqatWM92/AfZqyzqjCVFFJlcScG8ryqNtQacPuMqOMQJVWF8+ljDp3q7sy2Ro
5MBmNk7a4RBx5Q68MdHnDjm5vWedoKXwODKh3Ya3ICQfMSu6PM+DMkCqiYDLB+srqOvXvt5FENsN
C+69uOobrigpBjF7s/TnCqztE8myOPRlA9a0f6aj/h3Pmq64JrVwDkcrlC/NplOZ1algRkKDWh1E
H1ecsxcaFI9bhg1YId3zA5Iwt+E1Wdm+QPWi4mW0/9NktlOfdvKQg0v13wKQilBUlaKflW51jN2o
ASCKOqFI7fksvTmvzmRV65BtBaDIrYYfH9Me6cofgBJB2ttLZA7pTSa6XpCjnc6y9yKWr9hTu0P/
Icy8wCXW25hgH+iEZeX5tV0QguEyf+bR/Fh3i2vafECdacqSZF5xu/00AUc2u6RB6V5cg8+QIXLJ
AYxZUtej8e0CCC0EMuie0LxtBq9qiCYyg6xYZKmpF3OXNoC08Mekz0C5k+/uTvPGr8iYpHkG/pO5
qiIgDsPnnCsjgFZU67pxNVvMiz31KjbYWgZPc0t8pyzKUTHTFLY+UH9njqiTWNDFWSHiSIcVMivs
SEKwd8DH2mSpgPgLF7RBx7NTMC0Qsa6ridIfE+v5feRUhf1ujRMSEW0HOUPJd649HKcZIx9YWljw
ZMf4iRCQh6UQ9Vn0xwCOOBG9waOkstWUvLPK40vCq60Ka1OeLdGX+bLlbOh/GvOFaNzm2MPOCAUb
1VPlKwPC4Xm+amIf/YideJkw7sg3793qv6X/L9cA4x9iibGNhhkuI4b6gb4t9eDEvhuZTAVK0YJR
yX262MYdRNydrkN+uLveFsNw/nEKgaXtQorN1PoDVcCwDztNIkSzU0CnBQ6ouRNKiO3kCncGAfZ2
2O7oNvUtTzS8XuYORYSReJfS0WeT1gzFSqMVspcayJW49GmvUdkncug6D0TJddXUuIDX0TSlkVdH
YqOfxFwE5kaysQuAIJm9kOL5moxQX2bGDHIrdfxFJN+AMwygs8ab9h4xrFPDAfzdz+FMUdhHTdMH
yHsEAUl67sB0pUjN1aLav7PY1KgPHwEzbJK7xRC+ZH/Fanhz1M1AineUILYr26B2FZOmCcpW/r27
/GPMA1Y3fUG+kCc3o2fZ9LO4VGN1LQOhO5bmbQraeXi2j4tIBQlTqdo0Nwb1hUJ1RbiBzy4UH1CP
rWZwQPIg/qkz37Y5+ScXMfwkSqC+Hiy0zrDOECuIh/YVRP6NjOgm6CKYVUjE+O6f+GR6rTQYgB+9
LwjJVjdm0l4gkrHtnwXlzCNA8EXSj8ZltccSFKZGa06ZzGpzdMnXunMjnh5ORdeWFmEuzf8Ib8CC
YDj8BbhWVOVe6DNuGYo1xTj7xwVFfsOBTAhDoSsFn6XdMxIgF/t0p9JYbuS0Bv4jHZSIlo6PU9h2
k4ghcAekWXg5Q/9C8Ju1l4jg/RtF5HfXz+z8o0ac14jg+i07/FoPDwS/5zV5pV1T7hcCyRmWLxek
g2m3Czf3FM9VNhPvyib8PSUlEQfz3E1JKaArJ83hQjjZGm8eKj9igs+y2bHUCXF56wN9xs8zzek4
YY0862J+lWzOq17Z7Ezn9e7IPQKXE8az5YAP92QswsY0LsKC1df5fWK0pEN6boZjrmzW4T2FRAYR
prm0cMXnkKX2CMcCS4a2mhau6M0CI85TTr/w9toxL/lL6i7Qf1DfCzJElFZWgnHjls1I8XAZOxo9
kc1HJtcbhAJGLm9UAZjGRUtean1ptaSw2JBRv77TGFU1UT+4eavxsHj4uEnFu7XitkpAWZNuqq/1
gxnU3k2QaY4IMLIK73Y07eSamU6+lsc3z9H2GM2ZpP28BArdY+RtsOwEWGdrn1MC97/r9DdjAGH+
FrX1k2rx7R3hNX9fCip5lc3u/wsrMPAUMG2smFGuRU9Xqv2iosGmbQj9ElsLC2J/tv5I1RFOWqs+
1h+zRS2SApKwSuIwptoMwbxdFHDkgYKonUD8xNqJkFvV1lwueCvSYId/xzmRhaEVuh6acsyIY3et
60rElwXAQu00IPrbbw30my6cLpM1CNr/7NE7vYp0B/4tV7bIRgMQotImYxBzyQzyHtabnva9CbXA
v2ds4c1uV9qxKDSxxJ8BXfuJ8/xNI6NZupiv/u4LGw/p67U6Cma2iUknmlLcVSC47tmBfsGy6C+M
LsyHPhKzl5U6e25c10ZbZ2+WXya+jbhOYqvIVZEIinm6a6NqcY/TCfBuhx18f+rgKQr94xNwfCGc
YrUT/zXErMjyAbEberimwZT2jaTKbKRYmFMPumnflqqiUhvU7WsT0pSr1WEYY6pfNxmnhfHDbR0Q
7qhv6u/LnH4g7yZLcoMxzXFwnhICpJ3Q0m+KN2Z9f/m0dQljmAzMoBWZXOl6Jh4/0OUbXOUKTngk
4AdMlWxqxGP3H8kYxDTuO1TsibhIIyBhzkatbmydtZYNe3JtWvELj8XBmQigA248JgKMGWj9X3Kt
vs/T4Fgh1FgvkUXmXFxWrH90oqq9Yowqkvl79x/Tb1YX/63wpB5E9I52jqb5QPi0luTKR1FZne99
MxKTP3PzaIxPW1AIDlz0bVpF73NA9slQreiApm7OD0vS04/C1doiJdfjseUFce5ekg7B1J7XnDav
uRFO1cOeTF6qK7Yik6jfZ6xd0ySrJUKCib0otgwcWLehpd7jhANrlCeXwQKgcgDoiuWaFHSQ/0Xf
BP1O9t6gsE8Qr0azxxB3gzkKN9c3NBcaIISxIngDvs2vSVaNx3V79HzNNjZ5ju9whZKOeGDMpEo5
3zglYZpuFzwyMS7s9Tp8BGEz5ZH4BNrQK/V1KSk2CJfocOtmMtxNy1WNzctjYYFkcHb9FE0YVf8h
/Z907mCIdiV+0zzQeqgM/rLJRzvCcYHEdVsodO37UU/v5Dekfs/haLPJPduZ/e/9XwD4fwRoMFuE
RPPkPfIiWo+w/ktsTsmR6ZE+g6af07Q2Ii2QB4cEx5lYbzHYdhqJG2FFuAg9ElpEWgPpCfa1IsN4
y4pPr5vvck4dLsHyN7ZWcbPiiiwbyD941brwd28+PfWD9F8yFCDMzb95Mripaw/Qc4CqR6Q2SF6G
H+nIVWRoASbTes+a7ZO9T/iLffW9DDimvSFg9ROx9Xzf5jDTJPAfAQVswG1vP0Dw2zbnOQlNlcQf
ERMac5ShSkVy00WYwrxLjH7OAIMBkcFRLFF+5MyviIzu/rWCdPFELh+VAIcuqlNtR3h2pe0vvqoU
hD9P17D6PRb2B9jItJgIdEx1XiKiTJBoEgrDhv+n8FElUIpDjO37BlgtEYy3qRvz6sBTnAHISTgJ
kvGjWtZUVLgsqw1Lp0J5nfmgbUjwzMzcOq06Lo/tZf37vGQD2yy3ZGV9d62OXio9wlgwvrl5IQsL
IaENXJllT/pUM08jneZ9b5bXi4YqLGpmzl9mwDh6S50PlxFAEn3GmdOxPpF7XM4Y/1yIBf7SaFRg
zNSFp4+M2Z+oIkw7PwuJkmSk80lNtLG4XyGswbtVvNRZtAz+dDU0WX1i9eUK1U73ADp2mi/PmVnh
EVtJMlz42cbs/eJ3zq4JQJRt1t21jxrWDxKjAZjk7I3n+9yGrxXzC8mo4AJRrty+Wb/MshEBIota
h/uwQlcBwRTOTpKrM/oAbZIlyQCpCkTLokgUQxCDjDrABe08PVOG0g4PT2wzRCkiw0Grqa22CFQU
IVqOTX98JAWsC6ugow/pVyjhj+YQD1LIdtugiO3zIzdo/QQhMF4Gibxx43DoooT1sqPcA7MDIetD
HaljdGwKBgqFW8qzaQBFgl36zwj+3zXr8PXuRKvu3OddA/zq58RATtctPUPWsEuxbicZ+f6V6WhZ
MyrbxLZPNxQoNbqdf4LwxtJI0KWQ0lEq1pO3MP8/kPfUzJ84/elzMfPj7zL8ESAmCNc/C6Ws5Dxk
8y1Oiq/wTkaFxaTTixvjALvVJibJ3oOQSDmM2JSk5CZDRCtNk8219+YqpIdE+P1G9MaJyWcRzMYx
D/Cm7khPaUHXPfdyCEDgSZrySpNpYSzvDdqDJqx3vZpjqcMc3jkwMajbhx37rBRpJeA5R+YYPiZf
Eyx60bNCtdjUEYfYJdqpvDV0pm+HfJqw9kPIfp7VfAKmfegm15ZPcQ68sn4EnSjU63EufGocvwHT
k5kwpRgpAwqPIerECSmFwaoXa/Nxi2QP8vTnunhluVCngijpZrS5GyXPvDBro0chI7GkngW5cmrd
9xFpvtEDqsiaHqZllzfAenKS0wYyaQl/lvpDkkU3QUiBSa5Y7eyiMpxMs0z3U/KlHVJosrSoKHex
xz+qITZH9BLV6ykBGn65+D/08Fs79FxhpX/g8d8C6qNjBbkRI1Oy3FlUKPQisih7WVW5NfyCvGxI
ym+gbB40n/YYCA12VR/KNFYL+jkRn7IhFwCltfUZ5HH1FKC/xK8GqYK9L0f9AqwBl9UQPfDqbug3
a5osCGzjPe9M3yvnNU2Xu7g89nmcljz+QEWIdxaBjK26O2/W/yBUZfpnjHZWZNexSxZEi6WJTr+C
FIQfL/YmlUdQxwEkJRtztr6bfHLS1/schVKEDSHyeyT1qjWum7MENyBH0yv+40ZGqjRdZFFHn/x4
ji3c1bgiOUwMPm4lgVczzo6jrepwYkMcD/FD4i09r9yqAigyGoNkq9dx20cVufMMZ0VoVGtOH9B8
ygpARfLyJepNOk0FikWRQ3KXh745r2aVh/3qI7H79aBeLUapvQTsGCZtA86rgMdx+JInCr0KY/li
rNAWaeXMOFRhGAYZfPJ8D8rLHD1KlgG/fDjDLSKaYYvL16XC0JtJUSHVVYYQls7JYs3vkWw6mqzj
2rNVw3k4NnO2oeESmbLQacqHIPKBQdL7ZFL1oiB+lf7cOza4tcxU6kE0KIAylP+xuXaQQTmiEYSo
jqM/kLxOM7TfjbJlelnK8+JgGLXwRnNrTNMN36jlbwyL1XpDecIUuJqjwqcFFT59q8QHrJ+h8RUT
9ephTpZ4F4X2DVZtLb/5EsZmeDBKmL2bFGGRyXAqDabmoOmIuKNzJd/J51gebZO+iiEplcPiTK52
ukdVkBc0ZA4f08j9erT7BovdZeevhREeHF2lh4nrgWv9PwZEVrOAnylZo5coCNXmwr8G0kDJCtj7
DgK7xQvE+4zKj6JGPfKA94jeXumI9CWwcQfyyYg/nbfhpDQulJEgLU5FTlhkQCQF5Aevm0J6aQBz
2RMQhbu6mql68SVYEPK7QsDrvvqYQRcvPrFX5eNTKjs7LuX2nJYUKejoN9gJoOGEOaq9pwBp4gP6
HSYPlpjvth2CXjNm9arCG05CNsWWiKijJOFUXVaEka7APEuA//VtXFyKBOljfyn7kXhuBNVmVvff
OKbY+Q4S15ZIBPphNAvT1dysQedHaDdayupaS+pPZjM+9PuZw3JhpFYtGsvwGdyxA+hHaXjRzFiZ
7EM5ahm4rxo/MlU5cHwfSS7Edp+S9MdNS3EmFIVI9j4uXC4UjTOqeKZ9x21FKJ+xDEnVhsQ+Q/2b
ufhV/LzRXW3UOCib/+1AdiDs7tbPQqfLKbc26r7EfkdcbsdHksK+Eog0wxGg13KeiQ39odgtSQYC
rOOSvGL+FpxMM8YiyHE54KznXakzYNRGPhF+gVZf386TST8EeTmgF0yeRqYVV+hk4pqZet8gD5yS
CKA5LtpiwGwZoghlIJAx4U8X6zB1sfAvOvhZz+KRnV0aqByE75hQTJ6Ts/2eZAPwHuKEHgfaBI4d
UWXudduKO0GxRc02ZITEctnLjT7CkeIO4bNzFRJgyZW7suw1m3KQAA3ZdwLJYwPkXY+axb3emdQq
FpxClyir56CLEVTYOMpZxlyzvvoc/klpXUsZfJWuFtlcmflijjW45Dl0cSZIaxT8otA6T9NQJzB1
KJzjeFxrjpoQUgiua30nB/4koDJSj3HAsGZ/nfRkEMMNeJHPoh8G2Rd9bIUyZGzb/W/TEbQTvxlz
KMSGpDfdO/nbznUpigT9z+F5ckzCd0LoSbkVdIdNSa2YqOn0egOwZJYMQPQYJSgtMYcq20uARaLC
L9myAGwe5e5jyKUsbX5hUUo6q0VoAcuTOyim/a19XDpKZoX5JLixfeAuk6fWXk+vy3bFdiY9sz0Z
IdoEmBlSMQEzbbDtHZ5+vlhB2j0abTe+qPunVs5zTK6FTP0FdzCSCdXVpD01DRCtkeCU65HQFLEA
t5fuBel9f6eu0wKp9iXORDt8er2xVH91vJM/1WgVEtGRRKQFimMYDxeGc0dra8tTquWL0OqORpbL
MCMQwHsMJiYqakdEALvSgUQLBL/hYXLlZraYTLdFrLEZRlNjTMNOjlrnVeJlvfpDXTShDlsal7dr
nAcFlwdpLq+U7l+gefzxMzBo9ABX2hJcMViRd5fxMYXmwnwaqvulFy8/Sub2oMdxMrp1aUIHe0kM
8Uldl+FMbNeMX6zmBB2wOxbEd/3FIPmTBPpRWENM72yv5oHpXBNN0Ey2cH2rKMGpyO77UG8Bxp3y
Q+68Yl28VH+26alxjhoDINdOg6FU7FlF7W8EKYzoEimbOo1yvJWiUgAZVkSQYAGeztZMrrFzws3J
At0x2OSncmOctclW9ThlI5DmA/ZThda30WKTlEvGXUgppEXEY6QvudqdaJDb+zQbwcxcYAaV453P
+sOEcHgTeA0hi/G5f1q1BWoevAaD0COI18UGSMG9R88kmy4CArCAVIYOptjlOWyYcmZmoOXrlnys
S2OXLNL7UptRCRJC6N3Jxm5qvdwl8HLaBYfnDCbjQuk/h5DCP+KRo8xDixU3KMA1v/60nZvw+6RQ
7c0xsNgyTpsUnIfbsU/vMFOzFVkDNK53RHPq4JSqHKY28NV856xwKgBsR15w6sdM89vNk71RTTRk
DsnBTjKeqd7S+4OK3JaQuH8jxqJpa+WBHpCxa7NNo4ULvv78aGvlqzVeXmRTISEI7ZYXDkxxodU2
oSEXq8F6fdbSATYKleZcg3YgW+i0EaXomHx+y2JE7+pa9SkwyB2mKSPbh5wRPpZ2bE1wlyK8dLij
YQFxK+ufqk9fpY+aNboOdHe1nxpMHsUyRSWAvAXhjO+nPU8YlEs+J+YkqbUtiuWFFizZnhZw28oL
tNBDqDP/evJW3V+qxS6MdaLu7QeZw9iHxDtrus2MxuSZ1qZXvGe8KCIMklDTToDEhOT6qiU8jXPF
FVB2PiXHWx+J8/Mw2c+/pbx/HDEG0h+/8DYbIeSNtcnFJPkKDlJm9+lb+weFjc30KwHY7bnjKXP1
DoA1XEphzd77dhylpO+OuiNI0XgFr78Wdk1V+Q1giFV4GMpQGQJHLluPKRkamlWGc+9P05xNZ3LO
4vWFTQfeRqqH6a69G2cBwuMPUJlovXdgG5/PIrggS4b7lPEp83o5EuGNHi48Oqae1Ho2N6bt2Y3X
xgGdSndCs5b6JsbhjSe5moo0F+6xHIJpPxKl5G5Bad7irHuhIj85snuCuApnpJc/FSyDBv94eKRI
NtAQqvvrWDOkii18d4rQMPZWVCPUj9GPBZmdvWEQ5BhBPf0LbLR6Duv10eaH3XaH5Q+q5vrxkByq
1R/2emocsyzgDqdNwieQfKLn6/0KNkp2KA9ZpwFkLiLZ8FuTkGmywyfGeiTJM3PozlZn9hrMsPHd
vILd5RAz93rvAZom2mFqucouwMKAG+8Bqwib2aItXzV3ayUCSB+jwCBTRBW+udFN0oBuOht3bRGL
Cy0zLM1dT4/boNXm6Z6B3dKdZaGRj6CWuFaxkL02f5341uK8YJq/nckPhqOd+mQmr1Er7dLab+KE
HNUQzHRe+4666e3KisybwXK9GgiXUYagxi9wguGubQqhD4dVKkK2df+ZU2BA7nlghF+FOrGJGbuS
LWOyeW0maXK9137/wqc9Ri7mKUQAdtbKSTmHeILZ8ZMe1pfYiYCDKHdJ/Z58PP9yqCk4jkYzaQ9A
nqsS/5oqGk/FeDn++BAc0aRGSs33rV6/gglbe5J4EVFVjmy+tjekSIcePVZv6NEd4iyxi6S1AhOu
t59+FHxUv0gYK26vbssMbTklZvmcjb9aAdPTdBo4c6U9jNzx/WKtY8MtNtQ4Gv3ktMN9uJ6OaPsw
/1WdgtH3W8pZtoBMj8yN3LmZCWO78Q37hjmQgWiEwiTqlli1WFAjTR8MUhviMmAH7Ud4tXPGmXPf
quiWfI3WqhA/B7S82JmKbjmQUMiqXgoynbWfpXv+fHZtSl1R34n0zdoiHCFK+mOSyZqTLYID7cBM
zjjwqatRNYmdAArTZ8nGFb/WHbCfA+CkWXtuamDrfa1m11pDbzCkrlAvr5SiJbtyjArmcLvPKcbR
ZkZEcMANMx5DI60AsnI+ooucBRJa2hoaUfu9qOudqjapC5+GiDTT+aEkaWG8Vlcli3NtqWPykXh9
Q8eXc+3qu9szXjy5Ty8agxvEirNZeggnGhxKEwagzZ/p4Z54kszl0lSb/hbE6VbZtJnaSeXh6Vt8
A8wUXBo/WNi8nv2McFiPdvVS3A3oDJIMIOZeO5DmjTmq4pQ+dpAb9o2KszYdn3622GA6SuXfhMNu
Z86lKUXSCTaYkWzO7c5LjkAD9ByPtFHrD/JqDAcl2tgwm0HphBtbCDV12KY93g4bkfivZ3EoWMrP
Ql4KS/vObucQKaZ8RVk7TccYZdeLOsBN92EfT7baBtmn5FjJrbXDvX6hbXKDKInCqwsUs/ke24iv
23clfoniXgo47rRcfrdzb0G2BYIuU9AcxiB28x3X4a1mQ9bFl6/pLl/eIm/Tul4TseCfcAaTaxuX
0RXhkNDsx3WdM3BtedPnTudXGSQ0xxpddvaHUoNW5kTrP8n0qp2WrfOBhkIGUrH9jpQ2jDrimCMN
JELx4SjAgmcS4FeZiBAvBfE94IdA0QfsHLaFf2jlYh0v+8ORfrzxbwlue8tsA7kt7OPo3DhxPp1z
5Ru5CfRoplWDwzdK+CmiiXOD6UP4l50itgpfh52i3BDMw11sL+ptXU/ZCXhjonGHaYm9+D2nWwVU
SS2xF2lTmh9tFr6hAE9DLc3v68mezb2CeujQRsBNykgEp2gZxnSnG4WZa5UZ56cCHGOOQ+wzKNZX
L6mWceQA9FE6LmPlo1X7GcLCI0F9Uqdl+LoBCR8Lsf7a9Xv41VFymXhKZGxJZ5HB7eTF6I0KSlQY
gY/iSrdCDcIY5hzpXM7efaGWBO+Qskyb6um9e0ScKDGMAQhyenbGYef/5IkmW6IxK8gSAKqq5cG7
TzCvIOK74UH9TXfjGuE5snxLCjlaZsmYIM+ysVzkY2Oqq8vUgSWn8MPaqr/rEkVhJ+LHvcZWCGqA
h9eOvTmiDf2js0SYuC6Cvb1/lZ2ItXdsl+YvJNo2cVR2rDdhtKbzQmzYPFezKLB/lP40+IlKYdD+
8Zr5PzYey1oUtBgw5V3nBOr4mGBbSZ6sVg59reyleepZ1SzR4XblaKewyGKWp8zNezayzHxSLoFV
eTPiEdGWCLRmpQ1r+vmwa1yi78+Ll1ykrxbfXq6R/Xp+oSIR861Fp6Cre1UunTtf9O2DD/+YZPqh
X1HcuadHCvgUfjtEY7vwwvPo6peEn9aA+UqLb7q7RMirTXCiRpIiciUUW7p36Ri027u2O22Jkp4W
JTHZ+djokt1Pnr8EbFsxz3CloJHCS8M7LiY1TxuO+/5ekf2E2OWs6Ncu7keQFvNDJb7G0lzscGRH
OJY5IXjjr6lF6Hw/wM+QZL8eI43bEYRi0F+9hOM5q9XaxBKTf2Dkmi/BFCBPOjPJBKAN/Rr2pYWg
QbaOsKj5pMct0qGLsXsuKw4S+qUiqVDyxmE/4kJDlZHawRoedGU9RE2PqK/gRIzhvWs4zMrt4rFO
mSZMvaEIdjNuLx0iE7P6EjsT5YeYqzImSJUGIWMECjWlCeSqk/ua5VV+IQ6t06PMyafUyWxqlT0B
huzNpKE8EaXdlSgcL4WZBIBPUywxYu9fSmD3YrSOx9x4QvjFzW+oGDW3w6+3yMgKPk4x0fJRfbfX
D/M4PJLwXnyUaQGA1RuuqFgqVQECOQ5Xtf0b1rbT3FBMstCuMosCuxXzqHO61XLdpV4hhb6BvTFu
v/6b3JvVlhlyQhF2MJQtmC4o0j+bcTVHyiWTH90eIhlF7Yl0BEDFng1J+6w8EkhrmgfnCczjzu7U
CDp5OpWijFxDhsz/jHQa9FqWfbuD31oAMkv7z2NpkvCcrJxYJWT9i1uMD6asTuyDWRynFybR5hLp
WJGqGpaEbfzSGbgjL0rIMflbEkCo52hwDLHiWbCqj6OVH1lHALvJbIAkjlP4SfrLCkt70qYEieRf
r4wteaq6KcNz1qInluc2kcWq1VxCE56YXCu86FgBT7GuEtCX1Apa5P/S5BIoZMqXsiTMQbmk+iuQ
Q0M+IZjOxQxpWoKzM5K4QGHJ1589c7QRwKFKJeVrWE/r+ssXKruwgd01cDv7IT1DeRi37x4TRvu3
zUvp7UR5VnOVPs7H0oQWXB6N37vHN1o4efHDwq3irmFhrHaCvAsquZNQXfhmDm6yF13ApshMtA00
V8e/NPS2cNeMjc3CRM1vMSDQ5xcJFJ7dPZrheEHjoXYfLv5IwjpFaTyL2YJqOVNVTjvR/zqD/A1l
SR1xS9IRdjWFO2OarWrfO5eJu4ziRPFWbXOWqJkOu7eQNE7Nf3AcgKWplcGB2HDcO7O3TAZXVG97
ktMkxpMJZrA/cbWVlzPRHe8HLQU3eTogcfpdWfOwV4kGzcrmL48ML6sV5Cy6oyHqaoXvtyCmBz+x
PgHria0PByVyVVshylmAxMQ8uXwOuruAQkn2SU7cy16G6wZ8te+6qrZeRSFHVMJ7AiBSHG9DBHru
XQf/Pfk9/T1i3cCq4jKiGR3sohRdoYmKKh/Q8GpqYV7gP+5TgF89gEiYFoZan6rtKrbhjMjysx2+
NVTxTNmZ6reUnpQ44lTySOm4WnoGxZFW4IIiyyq3YcgF9ZU4TKZ/qVnieuoIVaqQyTOCTAt60w79
0bgQygC3Vl//Zjg/SPl70tHJAued23JW9/DJyTcHbkvOe5Tg7qrJbeyNeWiZDOhXLGaQv+L0fH6k
EwOwL6DFUxER0ruFgECUhTI/SADNh38A4fu8trml5Yl+wfUr2pI7r8cbTOcPFbPFPTHC/Mmhebxc
Ajhtdx6TgO5/NooJDNnrpTcZGhTsQZwQBFsIBhs/4/m/ye63WisXjUqIMRXX99Zvy1feWRLevA+W
UzjCB0hyiOQluBvjUtCGqlhIOGnYVcS79sUZPdvOpq8Aje5GuAbyMBdYtTiZybTh3qfnodrgKncY
SRkkUkqYXes2gEr+sMS3nU/+q4AWnzZQ3If5VkgfIwDZoxu09vDdUCQaUFwcQ0ZCJcEcvbq+8vTj
HE/fcO9UO3/+OCovAiOzAF9U5Ryqn5jGEVYVQOTyMmgXpuTTIjUyBA8PAWwp4kvjOIE7C/T+GcHs
32ght3X+/efNiQcIgs8f+sVeg2t2uFt13zj5Fx/74lN+P4N8MgIGSB7cEWh9hfKA4gBkrUR74ero
YiKWd0MOt+XJTrMzaM4zP1sp9k37Jx9Ja/LCB93DdWQ1lhcDnW46EOPsHzhVK6jy8vrsyf+QufrP
C+qwM0kpBr2CJFt5c9wOLHlg8ddT2LQnjLSyMsK7NjFz56H3IO+pXlQNPuylIyVmneM+quAUBzxT
FlIDoZXzJzN1nigI0RZtCaPCEXzJYZ6Djn9MPCvoD7XjInYsjsiy8kHGQHnEQeI7VETQuMHyLVCK
eLcfs85BU+uViPoUGdqd++QZsHAAlPHH/5tAsE2U/K3e6+aYh+snuPa9xZQOTEfuxi+X/2mumn1h
qiJfzVabSgXlXsMjPdSbeTp1NVxyXPYz0Nt9PSQ6KQTgyOXBxaEu+tZYq8C2Mds7iizRU7fhNQHD
MwpT5vaMJo/JMPatPT7sJA59sCLyLze0L2zlbRjJFEOfP4yWvaucFMAzkb06gD7bLQA3Vq6E3Pz+
f59tAU0Q1SuPJapM1Tk91+e6+U5KJhealu04p8DI/qZa6nNgseLewKksRmViuR6pY4JTjfLLS6M+
PDZbqLUjWQDUWN+rTIlxa+jJw6RmIRiqQsmOslJuPQeCtenpWEK3gyTRHUQqo52ThSDqULNel7s1
HNaTZomgG8CrNjkSlBwH5PAROli2YiVS36hGATNC+hKOHS4SpfWCp6g+AJVBJBtc2BhxDPo5lAqV
moQ2tTks7vuZ9MTrnAk/Wt5gIYrmv1kjwJSy5dFPrSjra4oKhmUBJUZrttGvlA5SGYxM2ogaUF2O
lfX4j/pQ+K9OwC/a080dcagOyx/X1CQna334ttJiNFYTH3VnyZOstQQS+sZaLjTrchDgfazvfVEu
r9CnrJisKpoTxwKVUEYazLXf4WxMQN6Tvy6P5Qj4yYGmlX2gvL0+xXOw2FmS43AjTWNyO8hOF4su
mOhtVU26CNUsOUUE8+HuhhOVxRyCbeOcAjSv2MYzlRTAll3Ci9W8fvJM2IqI0yx00OJqvj9PWfeB
+HhJSRMZE72jAyqvey6KMM1ewz9y/SuGJncMwEZV3rkRnHe7ElIOmSrF+1jEuSCnhusgH96Y5Xsu
qPHYIQcUsG7upUPy3JChUVLwZDK8mw6BJcdglVsIR4WRlGxCIAcx0w8M7K2rV5ZgAxC8jhyI6QEF
/v4VU34w8OGgBb0lIZz4ycwq7vfHuJrSCWKHwAKCjwrpf3qqVGQXovEnOahPjl6wUwzZoZodBzmK
te7DWGqdeFdKL/ksXsm6jjclpYYfQy/dE1k9ukUvOhkvc6rf3K/kxVmMxd4oiTcVSmpP3tQbiSZL
ZxyFQwc8ixT7U0i9hz8I/3clVjaDD37YrR1Z0AyT3l7MHg7q8cQF8DcrIuUzedNcZWvxypBRGxXZ
WVOX+9qM/wCDs5MBYRSAzTUpwZKQQJeynPatu8gyQ8qHR3XRdtwKFPbSuYfZ+2RMVrNOZppqDF/h
nWqvIm2hKNBWYX1JrDg7suW0Pju4bza4JBeWqFNrdkKIBJeMZkXP0VaGDOeROMA0JMCfTXe5Ynm6
aHyT4ICDiV3bQKw20mZUD3dzDkUAv4Kniskvo1hAs4vE0Vt7rQRJw+6S2jDDXhN78sSvn00P1FX/
mPv7/2Vv2GReoYl7DGOZF0XoVJVGApVZNJeakN2iACGQcStYkske95+nG9mftd5fe+u5UkWtpNLB
uZTTkdOiA9wP8axifKT6g/cvgFmvhKLtEPKkAiisQ8aIaQSdkZJCAD4s4CSxwbDvZVPjGZKndTlA
f4Aq/mmyBf9xTbhNE8DnTBkvAPOlIrLeJvfRTfl6Kl1eYaZEtWIITDYH3lfh0j4ypra1PVQONwBk
mza6fZz18GG4DVpT7Du3u5S7c477JepRoowQV8i8/M9qS0OeEJdvopL9VbBsqsB3F2Mdm7HcHQcJ
g1tTHqAX1zT/0F0Mserqd94KfDaI6qJnOPw9bEkOeHMT780FFn4ms8HzjP49MgJ2dNzifldK8FsO
FMSU4gj1KaP06aVK1mK+Z3+oXCP9NA26DQc/Y6ZR2n3R5HUz9VPAwJWsJUJ9T/FYNs1dmprndj2f
gs/tH5Y9Lvj2nnlwP6PSWdeSpkSAg0VVpQ6urlFgoR1cDhZfdxRBidgLfLlBYIWSHK+VVkNFS2mN
ISo4GKPm9LBfhzq0TmNmFyCCASLSLFy95TWLxPg7+KI6p5hPFZCiLrZeZ0yG0Nzr7EWcw/fB8Oc0
tRducVqOQCyxWsRzZpdWaFUSMPNwrrQt6FpjXBxytumL0FUg+cKqqQ2sJFAS/5tNLizGBhntFfJX
UD5A1BDdHRd5nXyehbKZcV3u7NxpiV6HdeIzS/obJ/29l/0Z+l/ixYz3YjCdxFueFPPmOkjdrI+4
PW1mCe5sTuQKNhFzmUUrKO1oDU2WeiavqUlZma5MIiSz8Ae8/haQf/N7tCOneCbUQxN16eFShr3d
YGAnI7awcoyst4W9iV747vYIGjmW6Th3MKFgOHARnDCTPfl+V34g27cxV2kPCHCOVu3xT5QC+lEl
4hgnbr7s1tGAeeeyFOW1GjoxRUhgv+4o0JA/OfMo7Is5nhOqTXZUmC0lp14VsjHglo5ksZxG/O9F
nEmHqRNUaVV39NECGz4YK7/qVuUtQ7W6kTKqWFW57BNi6GKSyIxLDjnJ6D4B/mZ5zaCz4tpSX2qx
jHHS32OZtan1dAZ9M3ERdhnla1yI6nQt5WB+4OuaeIxBnYqJi73rQ3mgdVVaLPR0iwpDVIdj4DVO
b3SA/fOpE0Nx3qdv9h6onVXWz59WGZv6jvZ7kATrrfiAJHYhDereZ4cf4WRc6C8VyIlNMpqyY2y+
XFk4hMs/Z7py18v07LD2QjZYiU1J9EAIp5HGVSBwsDzFfyhfqyi6nLs36ei+n5OgtXoNXkHn59mv
BwJhvaYuLb6CM5scPvnp2x/CXZ6zYLkx5jYKCdS/cgAjsY3L/d4Pp9KQiPhGt7fwv0+v4xt4IdlT
LPXv8BWsNU0a+zXLgmBErGd/futXByUJ+xa5aVHwuctIeS10u27hV7XBGfwGW4X8tDsDPbtxgv2/
R6cqn/PyjYWWmQx5Y5VZMqvRfOhnXHUe6gfSrprFc2rPVn0ny/i84MSz9ej0D139ystf6HJD5LIc
lsUUaTSeulswK/JNrlZYHcbtykqFYyU89l96phmo/FsXeoYhIgsOkRqT97wDJKv9pmID0q+2cGaK
qglIjkRvL9QoeuyF1nDG63D68hk3kVR7hgZPoAXf1NeIKKT8lLmWiPVILI9b7nzVNFQp/jkj/25v
al0yCAbsYnewWWUpw7HDOEjjqlW2Q4zpnF4p5rpUHEPb9Pc900y/bb2PJRlOv7YaMIyQQCg9mKud
pYSbHOPCmKpNsZhN5G+2Q5z/fXWa6bGyea2SmJxNdFVW7NmOvfnha999TlNiOLZNPzd7yZkbDSVf
aEhNQ16nbzv0W5D3YuplQXAcWtDjD0QDIC486Fs5lQ/VMJIuB6RBCB+Dv8SAg0niSkTaHwVSGOvX
njcbMjV6sdRQRbJJzIg3RgSOWEgAl+l+VyWGkeRyC+ht21tvzgjcleIEM+JQmNZi1CHmUDrlPvWE
Ibh5mYLHnKgqjAEdznAe9tc3cNrS2piXUgKxCSk3kMqiOB+/1wLUQASOFaUlaemY92XjJCo9XxUD
Uit66nZfgNv313/PoZoGcR/mwjtckwN70FC9UuYUzSrn6o9xzOfnO2KSd2QwIX3kxyCQC+syOPD4
jW6BHH77kLJX+XwHh+KBpaIP7yQE6SBSKRIW4vlrR42ckaQQW1RHmG8JAzFDl0B+5zaz/XPo8lNQ
I7rX2ic4Ac4Zg7tLwmkpFYVhF8r1TPBBFiMO2Lnll45boSDRnaoJbQ8PddHGp89SS6mohXwUla+i
Hfw42fW8tkC0ATJK3cDqfQI3wRzWvObdmdfFLvlSNOJfPdiK1d3naNY08oSCDkIRFf9+S+9z2E7P
cPN4oZulXMEmo2EvxjCnV858Idv2j55giaoLREUMTrRtj3ZexXY5pjpMaqGoKsRS+1wvPqiT48J8
kS6iJXI2h6/qaZGqWk2LPX49f+Vwp5ZCCetUDdlef4msIAV4AxyhMv0X5sBPPYtCB6zLweXEftbF
T+CmvOHNJtRnqZRlIgdsIdP0sOrMUzmO84LygsotlibGTvaHk+u6I66HwhS0TjZ8Fz3wbzlsIFd3
mYprmXsGzmUbooCCmkIfDbihOUgbHI48isXrPlEdvVBO7RUiHu0GtnfWZebRxVrSKlmM4Yo82YwF
nGZ2vZnk6nIfHRZBwpu89h+j6FAld7RvldZvnTlVSGGHbUeO+933OUfqT0jUJGOVQlYWl5jPTOCw
OJt/u44TAgTE7xpal2wOQIGtnPHX4PH9KbFu+/5zuiN3LGJ4MUeIyf9tbxnivPghS+L2J3tMkRz/
cOYz2PU1+1ExwYuuhsRebjSahOX6N07WU+axgz4mTzp7lrVvGg9bXU/yuJkUG3fS0Gh5ekAn/55I
kctdxG9KOun38rKCX+RsPmzOpoGgSqQH5DbreABI4K9EBIbAq1avT4Jt4ZFRd142jQOzRtR6yKIN
uDp/NAg8xFhZMFTyRh70vR8IwhhNj3kPphv0VAnCGwDZsin49DswoHlMU5v9IjjAkYZV8pqzygON
GJzChyXWLJaNzShDGeppuA9MTnMiQYz0hNZLzUKTWMu5fwtYISScCjqwEBCZ1YCPZ/dXS1DceCAJ
2Dyo/R35yYY0vBTFbzhaqBO2GqcLpaF+HshqFaN1Zj9DEPMs28Gd0oQodRUxGEKoOfhf+r6T4RT8
DnDezStjuTr1kcpkh9YsYRr1C/k3qALXv186mRqqseQpXUXnBEwx80fA/Sh+2Durd4Ftl+PSWoSI
nrn5YZA5fkg2gP5s3sn52ysmM9R5tpkHMiaAdWPcVXazz5tqILRr6WpXD8L9KBrfgW+U9PFAV7KD
a/CAwj5yhht+6XCYW8CpMIlyj65O9whD1MNNNcHLCxemloD97FwYmm8l6OiilggsHDeKpeYOu4/0
GAa9Me+zbZbsoZJcAfbtpW0gc/VyTpptrIYCw7bHDkChKvG9NyGQorQJKbX7GUMw7VothNlRrACT
X7G260MRK2Xv6EwpQ6jOB9T7D9haXCpNyTxCQDFyGceLYaxMkXA6m00irJPqQSoBmbVy5MQKu/LX
qU4N5dtbmo9c/GHv7Fbb63pYxBQAb5Y7HOr6UkhShiNC+L+233sZIH/QXObEJ63VnTUKKfyG7q/M
ehEqVlSbaEpW/x23RfM3GAX40joG4UDjhae6TqUofqyms+t3SE2EbEaO35HsHfJCtf6VuhB7lvMx
olNl58Bel0LECn0RpbOh4EpYLlv6iJz2iqBNBCm89LYPysqbxG9KLG/1VjpvwKJ/pIe8HfSYVMfg
R4NSoxuBPG2fn5msbdvjo+An0ck8z+mMwcf+OyZ2VqS3Uh/CAtZDeQ1oAEtQA5OJ5/7rf24QRcpf
SkYjvOxrqTVYe1ngxeuUyiiC+h0OG3p07d1RTJh7mxMwMt/7aygfhzx/sG3vUW/ph+xJ0Lp1aimh
Qc1tulR+bznLBcLN5Hc4a8xXgjN3tWr35uFpiRY8T3wPfh+afxghA8gLEsvvNoaHq0JAaRyRljyF
5Hmu5Tr23V4pMGHr83LpISVOA8zXNfjePDooon0tt5t/hFr/q1B+PGRbXc1whptqFibkLRmEyPZh
V3a3gHqWm1THokFrZEzbw4kcR/VATAY1bSAKBLfky/F0wgibYDMQgXhy6bBfnkDpnQYtLFtl+7u1
NJiyTDs9Ue4l/GNaXI9MxLvktaLVvJTxy0rcMZW68AS+Whllo1M16d8VaNxNRFF1QfFBvfkNx9Hr
eJJIk82oJP5BHTxvWwoeOzH3CUmeLW+OnB/8gsZCPCyPlJYai5WDNNbEYo2pf47uLUjLO90kBWkg
WnwiOa64sgsaHg1YcoC7Q+ZY+MGIgPE+VbHs7PdqlERA7a2xNmCkZ/3/EoQsr3lJE/Y47SDTT0Y9
cn4Hmq9w3gS9DlR5vbksO/VYGLSf8uvmOrUaTpI4E4Tiqjm/bbDSbV32aYREAoq+4Eg6TN3kNe4R
WvV3jAE2fjQXmfjPi3MF6sDkLAXj4+g9XLxSXizmSgi+5YN/o/cJhKwokWcb4wZjgwa78u+hLlMZ
dQmzC5o+08S0Ps80zXcxgQPgIstRa8daftPOZ5z8SmPDiSnG4V1gA7NXJCbNfOeBc7on8xIDievr
TXzP3l1yilCDUDZE0XAQK1VXMlp7LhXbKj/CbN3AydCimbkJhZX6thrpbtJAwMio0ddDc5UZ+F9z
NIPHa+YSBb+Zcyn6nCfjq+8v/k+eAilmJtp0sHGlpMXIsRqmqxG/RNzBad8jbi5k3fLqXKwjWFjG
ken1gMERZx+0FK6/nx0CFo3fFYa5KUT+luVYU1pr3v0LvYcIRT/m6DX70IwkV7JU9Fo6UVRLJzmM
OTwF0R2wr8Xkw73aLnWggwCE/q+nq0TldLS/Y+XhntGhVD89ATI6gLmFSN6OA4XfDzTtjZg5dcK6
5nkqUZEp/+2cGKn0beXCpNhzrosep7lzTo0LxlKMM5MkC6kOrPEQQQXEy7SAjdfLS+H0GHs/mjoQ
ocM9iVKslv3KYk7bUyEEORFr7TjWmKNTzQCGHa7IXbWSeAkk8BMOx0L5yqwFWbxDZIY4HlnsDxLG
OUZJkeTfszFSWOE0+wTvSIuVua2BT9PxGpBtYAS9vTQ4nyquXJTZkZDUhYY/ZqCoBh3CPuoM+62n
ZeSMf6x04o14A2kRW2dh1kAxnr5ear+nxt9a7Rdb1t75aOiFE0FaG+jq+Lbd5mStPIDnZn8TOeiv
E9/sW5Vsim3WT2+V1eKYqvA8fplngYF6akp0pNBCqdKm5ZTShfHup20DO83i9XySSGQ2yhT8EI20
kkuhlNr0KeIASoiegrQBf1ySE5ka8OnbbyscC8EAVnsQHQkyIdEP/4QplY9JRzu5VdFus0t2FdV7
HkJa69fWgEN9cE/OIE87KDtJe3RXGQCsh4sF7llqyEWjRo7LgVzTt0I6sVJGQYw34wyMp0oIR3qS
z6VDdmNP80a+ZMN/lf1ec6GVeSluILEq+oRO6q8WugCb2LmDK6i7m9WLl5/imayzH4TJXZ9K1apU
c+RVxPiLC8V12VhV4NNyuvgAIkwz5cGFr2jqdY86EmkPDWaoL6nsngIiYS6WHEFALUI5wtT00aHM
nrKJNNCGrNOBC3sPKaRY0tOydzRW/S0JQ/HxZCC39dIJjL0Jv63Yle6Dju9GQBjS/8obyHei14IA
iOnFjxMbJ0D4KExbffibfzCS7XT/HCKGjWWjKcu5t3Sknu+Zk8iSweO2e7Xf6AwdjLLOoxUF+Yxs
RrlmzriXtF82pxoEfEk1hqHI+2KAA5YL5FQBDz7Da2PiNPQy06bhYqmvumsNeU9Gx+zXKGZFaoo+
I+2NVes2xr2dUQKfoBy/BHzDznF+CXpWRwlPW7ommgPFlPYHPDMxfGVuBAPQR2lcwSZ9d4xt1SRO
yUITq+Uu8/BH/Q6MjIYUg2GxAnzbioU4r3pJxnZG6fNhEMHNQ7BkDE7LXYPe3dOFck3Of01nP0P9
M0mv3cFF3c9MLwSFbaV5JQ+LAVj2C7YjkQPW31ra6V/k/IHwwwn/JCLpCW2m2Ich0MHMaCIAjGDz
DSw92D7enny/t0/plp+ea4O4t5K0C+FOZl6tVmkfNeCdI8WRuMSlsOMb9PtmDFA/2GtCY//qXMUg
lVFRgOucprev5i7/2X0xtYMsZRahwX8AZH1SzXYF+szCbV6KsKwhqrF6bo4kl9AcEJliUf4mgxC6
CMG411zzqSmIsnSKNRI6GbxuDciYYcySCEpcCpTMxMaKHCS+oa0J8RkVXGLtiMsd4R5SjHFmhrbt
IFHNAe9MHvKjNjivJPbMO0SP085UmpGnIdDoPyddYstBch5zhrf3E25RvJLkM3GnsHoDitO4vR9q
9vjU+w0Ut5WJzR832ay161oMDEJG12PuHcLnfLTGmq4zIbDREkQGK2ScyO5FlC7dNop7wFPAXClY
SsgbwQv4awCObxCp3VLChlyl73vauw8vkazK1SvdY2X/z2RnIdPEjFbZn3GnZBkcRLwaJLQo7nNA
qPcxXn6I+rf6NzD/seTyi2hiN6zPOZH2ZtvTGbuWIsoURpf9Ayi7XvPJvU9ZHlAV3YjVS3Za+9KZ
V7aT3EePe9WnYKC2SjW2+gUagRjMkbEa+7Gcg+yr6dFekfV817Bs54u2PK6scVzGpx60oKSTMq5V
YSmPMq0Nhl3cz1j6QTNiX5cMhjeCfaEXEHBFzHj1PNJgqCVtUWzazoAnR3YYPSRxys2Tjwu4jBJc
EHLuUbcHM8kvUa/MZiwwdJk50NDxMys4Z3CSWoAGKxI45EummMjrouxSgS79h6J022a1aHgg23fs
+6jq/kokixUycWfN20X4l0kf5m5bl6lZEd9ks1uJzyBpup/yjorRQ+aYuFzO7NfIPqOyFKVjPTZ+
DMY+8RRiso2N29v/7/rd6yGvJxAbEJLhvQCYWy27hnFhJoEzTiS5+AZAK770ANIoq7jatHGpm4S4
Z4KGylES+lZRrC+snHMCgwe1XMs+b3nlW4MqeoQAzTENIU6oE7vnfH7S9mj+pzIay16bypOEEmuV
N4tEyxtRw9ywPRmKZlZ57N9tdRzh4CKu53wzErGKTKRsIaIzM/hRvd9CsYpuEV1M529cK0ZgbuRH
tA6JiOCLZ1Xy8JIjGemS7xmIICqEOs8mOgXFAY8tflaX1vdv1R2+smvnqJSaNkPfSTIvOSZ0L2hZ
S7V78YFyhcAYNU5LeimZVx1wpbJDp3omacLJqRWOREBMaIaowIzjLDehiSoDajvhMNy5LtDWKcvG
97HiuQ1G06EAg6fQs5ZbwN+PveUOzKhsX7EdZBMwCxZm8rZXUu6yprbZTHNuQ9vkCPcxtebWJv4f
4KSZrv97QYmpjDMiH6EnnNoka10vYfJekbplx5UDBjTT7fU5PSID063zrObRA9HTAb06plvLr5X9
pPqGi/6WHgJ5C0s7JAGbPnU6av1AJe4aBXcNb4UY9KjfXw8cOY4jdWa9wnrIySrrZgWGOG4uSeDb
fuB1jDMXu9YiCKFi7Q9Ynj4Wd/LgCy4X2i3I23AfVgZS9uLo64iSOnvDy3T8OYDidxM+5GsSAHzM
6Il22cFaPMQtnlx4HMqGvOa1EEUNVEF0+rTK+JE+iM8hEzVvGJGoLmxOdXEnRgivahHrVqvty0Br
eP8h3w4RwOLxkdt6rGcbsaFExrykM2CDwJSuh0x7635k1mTN3XwRn2/KB7XLa2A3dlf553cFPVnK
Ej00TSoOW4zReQnSB3iZ0Yk1bNkuHJd4xoZ0V9kn7aCNVDs4c00SiSVD7N2FG8xqzt4l0jjXtxmr
mvHxvrZt5DcXzXnCn/SFeF+R1TbpYPYfk9/OhZCg25CPMc2WS1gWtauUQ2SaNG9s4qIohjhSE7+n
r/7CyoM/57BCS6APj6hLLgmEcxnty3MxoLXS+gLHVy7xl5bWqNRovfv414jOXjnPB5Z+BFCQEsoB
BIwS0x6GNXo19CkiCJVUEFtabJQ+3vMufWAN7kmwU7JSqlky0qVhZvTHWk3eatx96mpsqI/Cp7Xn
K/dveu+rJB42WzCNI24aa6p316eo0VGgaMpNHQ8tD03DGbCweYzLL5lTJA6cC0EU+waGqIXbz6Gk
K+G8pr6d5x9ZIjrkRfsdjDBR40gZwvEeCAQk3X8zgiPsV0JknhU7JkPCn6zy4AmAa1h9dvBT9cNa
Zowb6KGfPNfyBZvjOAtt+j5ODsOqZUa4g59PiiodlypWKFpzcZwEq5FcxQodCjdcSs7ntkZuxVOC
eLqAJdQh2KM2DNlgCGPcMn6mg9gQBAhSd/ghTapt76LTtB8ve4Gb0NyhxoN47bI9HGL1/OOUjLiq
hCKPgB4/2/QvhU8JSqsHztjqFJbPMbGDAlJaVhGfFiE8Lo9At1P+LgA7ro63BkUjritnhkEl50+q
jt3k9UfPj9o3piOveGr5gK3gnIJu8E/CkNlAw4uWA1uMqdtgLJJptdY4FeCkEoM/WIYDi3f++ELO
xPAWksnqsl9Mzg28ubWFlqGWYNaoHSscEP/UL71nexI7K57PNrgF5JRJEatwhBSJZ/1sOncT3iw6
JnX7uIckMFCoqY8k9RwXxcl5fNmAvVj0+CY5RldoNk+EB16i0HtYeJ1V05jeJ82TP5m22NhmWiiq
Ix1Kxt2EdmI2tFTDGOs6QakYpfbC5Qh/faSbXWRnme+qBgc79FjUv/UrdXMI1P31V27T1u4WfmR9
x7f0wvf+mXpb6k1/nwCTgmTIUbOmK+45tqLojZ90diz5COCnZaviQz0H7camWI9q3Xye1td0jq+9
FBByeTbvojg6bQ69BmUDfsTYIb1DQKPbwl7mzJYeggtDQrLxKzGYwH5a622Df1l8Em8LOa0pqR9y
eTz3aV4rP01nx/5C5ohr/o67qQRlHQ3HBaUVkjJpIWYBcbJ2A/daodhAIKlMpaFvfuK1Sm/MSJMW
0Fwr6R4Iei4XkkH0kPGPLBOIwI6qaqfqnD6yJMsBuqAgqBsZwa7ibQ8/zL1xvo/QKjRpEA/BVpjH
i7OPQoDnFX8vKPYfq/hIkpplbYZKKmdpU7UOqf6ullmFFSlvdg9c01wR5jPFKVisK7gTwR+2jFbz
FWFy0hpfqZ6t0nsZfyLPrFpg9gp06dE7On9qfY8orGmun55vtVTfKzXCqPVor/SAfjBSWI9PpEr4
qZAsFUtwopwS+iatI6AZ891H4zJpzOWlXGDy6iTlRDumG1BM7ngYNByr9uhXkN7j7TaM4vqLckwv
T4fJSI0EZvB8+1ow7CtfRkRDGa+J4h3LBV+C/aJhnK/K9lsWA+g3Scj0IAA+ukA3buAIxxSzMpgD
A6Dcb8FAk3HyYrr0/+emJiMXlOq9T7h+R1XCD3ThnlPZAlisD9Evg/HIA6AXzDiYz2gbJJdBvkWJ
DWpaZp2D2FsJxq5H/laBiu5Tc0Gus7PyiJmaBA3C4LByhp7GzTuFgmjJgDyNQwyaOaU9UNbYWi67
M1FBayoFTlUTt6LM1VaKZbIKsy00BRR0DArxFWK7reVZkq9GbfzohrS8hoQ8FgQN7hzKR2DBNIdy
zyYCFYb/rr77NJd6TIOxQM2PF/mAEUOe9Kq96yHcEy9JSu7iRja7VQ8JVzplgN+hO8dbCFcmJ0tk
MdPYaV8iuzsZ26+xxk8vAG44pf/TeMwIY71YVROQuctQaEvOVAJrGu2kyrn7r21ZiL542aHcXBTM
tVLptlvFbYyxbOvCOg4/9aymMl8okfW8uKevdcvekJDfZxR7bxxHJZiMoASiFCuHcZS0u9psWunC
7+fyYpRawCk5C81cDG/DsnPXUck+3PemiovsLnWkGFphdR4Iz+Dob8kXJ6PUhf2UHQujVK0D///E
6QVSvdk8/y63rQKdqkn7rSJv69BbTToFIo9zv7cuf/Te0bYFc6EzLbUkLdoVb+LGSVA819lb9ozI
ZMfsgdEjJZg/jl+OlbvSEHrcff7mPj51hC/fhVrlK5OLbNolDxvnv7Ru1GYjjqD3F76DCsHlclZ3
gVo5fWhuRCpyzMHFPM9eeWbmWszqkM6zEbmmghsJskHp0YKWaaHw8Bi4noTi5i0GYt3co6SMW9zX
mDC9S3pxdlQwtiPecmn2Eu4Sp+LheuInCv26zs9iayGLOLHictuTD3ZYKvtTlSheNQhEBwZ7YHYv
ZKg8qKsxTvgBFm7I3K+4bNGIRTrguZ8o/OtUlo+ObrvugpA1e1cdXodClVwYCZQoFg/Ia9qEjwsY
uFBigTBSCPJ9E6e3uhDmStJ7G1+KKe1awB1RpvfJzspLRBFpWfVb4M5oXwy7v9YXAldjluXCDSXp
YodkoVxoQAvrAEchQOrXaqIYkCnRamvmYVEJgk75OMaNOZBeZ7tdnhzBNvEgOC7lzwy0F28sHJgN
I4vcSFjzG/JHKhrlvDrqYEelssKKyBOQFmUYf0rH36GlYHWLS5ejI1ZGs+T9Y65R3WmlS9wSv0eR
RGSwkkuMfBWHCai+xTvSUudrQFndmcfxM58lgdyPiwQBhP+eCE0YwIaxr3BIipQBENUxWNnG1xDb
4uEBbv8mRYnwSSr4s6sYQyrNMfkYwYNTnkYA1MlKjsKLpi6QnKGXfVfQukafHt1CE4ZBA8SF+Re3
IviCBPgnrGuY8HjtXVB7jpyLm6Bmacif+Oux6ccHGlf06i7fVQvNux3Sb0p9JAjbD+6UYZz9u9Je
WYfIl3CxwhHlDYR6yXn4B9liqNwVYinH3DanoDO4DwUjKE6JBQpUupg4FiEq2AGU5FAgES514Sy+
5aw2ml+Xl/9HgB/bSxQSVrVVuDs+m26Gf3KilF+g421DxETmESs61RgxG3bK806njHS7xJ1TFVDE
vSrhX/ZOTTEoD5BV/IfTBwdovYYnTe8320bTtFaIf8kMy3fsAGbH3G6WySYP/vDeFPlsJ47T968U
Mm0qtX39DckWUIIt+bOQLny4iy2j5a2MHhoSqqQvvX3aw9/RzdufDyTN98hL7DcmlD+/chR02l12
X1/o45UbBNJ9nXbOPzh7DDbCX0ZrgsKgOxec0T4aHEJbFMPncKprgx78MtUF/g/poLx3gMfwG5dp
ichh88ylSfZNYQz4ItGuYuRyw3y13JW65xXb5CkQtM4WKxCRW56zKE/aQr/wZKEUqNCIOH9UNt1N
jVpjo+H2PJmPMqFjnk8AioNd8Dj7bY8pDSVLc2uqfOsDCneLaKWMfLM2KihBGgL5MaaLlSHJLuQ9
S8+4RNPxl4NZjgP1nPkB/0z2iSDPbW2qnc643DSomGkShdOPLFc9k1+zy86YPw1PT01yAAl9MB81
YiJHHnD3ulB6OmDjY0YIA60DQ1/Kh9iRsbhy9bzn/4QbF+7zfLAGFuo4A9C5954SGhk78hnYCMa1
XGNYFYWwDLNkYQbcmf0zgoFFyqCOYEm2WAbhGFpHBmlsVhuBp6vcxolWNvCTIJcg8+I623Z0obSF
ssZlk9hlCEeNiniqTfHLv4sVX3hbPNF/8KHJtgvWEYjh3Vr+W6Z6faHiomcCpj1CPGO2uDKNB+CM
RBfeJYcpkl1V/R1k6WEsZhG5VEfMTv0kNTt83uG41gj902AOx4s24r5mMJMNjycj4PVrgOn3bRhJ
pkMYFKGeMzsKMfVO4nOGKSsgxFdSJZAU4OES8jt/giWmKP4JzVsHCjQrcg2oeb4ncF4PCs8GNMv6
MZwnGg6esngxtH5clBfzAWE91NBhX+TQV424UErSakX836RGsCODHX6qfxxFW1vAmZQI+WfdbqFW
zQg7FNB4szqDd0XLMH3nHyDRDxpMMNdIF/hWQX3qb4DnT3DOk/exRFMfAeOL4UUjtuMDGAHtcvBD
TZsd1u9JxIY9PpSmlahYQusFBRfJJ0IAvkfIClL2enKmLwTgt/MiyyYr5E5TSbhFUjxkC/NixqOK
mO0utm0ksnukyJWgmUitMql63IwWqav84dw09yKHJO1m/VKTkgaHhHQqj0AQBR2zD1vWahRxh+je
Vz0gRlhTGbYyXWpJH0fudGOd8jYF4PEDIE/BwHfzZd8PbF54PtJjzeMCcTBH6NFaL5u1+cyqyLu/
QpmcSo8S7vsPjcxv/W3MZTZZx3XTgVFzBAXi8THEx1BDLJHIXjPnYJQmkemH7aZz4OyLuAQf1EyF
SipXIB+Vf6U23C0TFiER3AhTTlVuASz5Qe2llZ7h4c5UGsqSub3U6AjvZdjrltZVEjcGDAr7JaQn
anfOLgEeKKsX3pL8XslzumTze2TR2J44DwBTe4+ZyZpaRoX1ZxMReUf9i4iSRANGW0jMfU9nxXxc
KgJ/0cEGYdIhB86t4/jGbkI+kEcOkMsrRGU+Bij0sNCejMi6xSr7OMWa80nuoOA8fnEfo9JPQQeV
3ddBo7uwx1FMzWSRRPXFaoCA2uffpRokOIMknIs9AftMii5eo8nIfz7qAkBMOu3WM+0+1tkGKL1w
4DAMTSKPj477o0kkxFJPDk9ykz6Derdwy4YEdhNaojdXd6To0awyrSv8kHp3S7IXanSPDi9SMVt1
P1qx/WAv2Jy3uS2IEViva+vSOubfFSgY0GkdXgO7MQPc21oqk8uvojmJGQi5fV1PmO9FQu9kXWHh
SUKMmPs+WZWiLXxbzfP7rwpQHWiIamLF3n3qTb+wNkjuZHbhDt1V1CY08I0sgROJrEDgNR1pwd/C
jBB+XJ3Ds6yT3k74W4QL/tvQOn9GJCtytKNKygHqMBcIPGAPArHc7oGHj4xag1w2TJgdQjHItQCI
axpfNO3NeJHLhKnX+PIOOu/+GUcnNkqHsvC0VwoVol7gwnkBXsr4DfDdw4WgeK7KdseTcg+lH+fE
UMTBOzhiDGR0zvFd4WAHaQ0ZApRQshMF9XRRS6H0metj3X6Wc2t2fA0UxZQjigV8iCeICNlVapIs
aXxBeRlLCS4DXA+d8w0rc4wIbqZU6EcRZ5H/TmF7Amn1fO8mrsHjsTpiUXVZw1qBcMsZuTyBWIqM
K5OIcTsnXWxN63KYT8w/CZSXmunfCU0TPdsh2dV7SQEO+1hswG/dZwze+cHZVQcZwrTm/1TYUd7p
lMloNBLVvz/2252qOzwS1HmKg/p6isgZzTMKfOuIk9OuELl9OSn1Zbm5y4F5E8tgBNvSc+DyHF3l
oKHKwmFZm5HsNIPF7z+cciJW6OuNU/fm+fLH4bdyYoX+ywGw9fngkR28egVqqWYjBWYITBBg5B9N
d9Cit+R3sKycyJiADbBBvRhDIdSBlWB5UMrPGNrdygU1YAC3LUHgzJmRKYeIpmUiHAycsDFgX80v
wcOHuHj2XjJsWsPgX03vkrxQzGHcOALHrjGS0bSgROh+Q/mhk8J2h/Ib3JvD7fyRzxf0ZXWPWXT/
WF6x2gPiUP9QhE3W8b7EDKF3h0Cn1rVndVA5yMTkHD8eUECvF2mMzCW74Zc45iYoBJIM+aNIVKI9
1wMuJqB6/3xfWcmWSOYiR5jCZEO0D7NosJ3T6Iohs0VktPiDhAAWBgTIOfUS6qcNxKGXl5mdX4ff
YHwSQv9ytw0mI8vh5x+0eFcSrbtebYuiHgIAlSYaEP2+YoBfKoEW0W8EQa4sXTkxlwvyxYVM+bt2
HzuyqGB+Pzt13nL+6QItiu4iJMYOKSFyJcNcG+XanPa/6HDpMxXcOUUqGFIuYwsi5/9fsrpE0L09
K9Wu9f5vfLtNwKc3aCtqUo3JR8GOAWJM43ajBHePBIIsz0akcxy4geI74GMU47TV4ahMKSyyIo1k
1SYMX5myOm04jShUYwsb4JoY7QFF1MpUuP/l4/27EZiUoHdVcvsezI7umusXBVPiVvnPZ5zXraGu
DDk0h8pT1QCPq3wghGvISbnTQd2Hsrw95ui4O0+YIfe4n3o9sxCSX39gzO3mw9CT9buAOHZDB73U
pXMLX9AoweSZP32dYgDhMse7S6sB2PGbeZP44f4JEJdP86OksR6K149DpZkp0vG2ObOHUYKLIEt6
xQwm1zx9wHQcw/d+nRFu0m+qzTh6m0mchscmUNXR3QqoTN0DFghhx2mHFMYANlyaFbYwSSpq8Smb
1CCWCZmJGUscnSyYx+k5i0s3DMsu6LnAIQlqUNwqdsr8FxlotK1iP3BQmdCvot7UeoH12aT2J6l6
Esai5ugaMk1tvtfJSIiE2Vrcbe/yoILYZ28K53SsFOxDw4zN5LwdroMlsnkusFxUZCtsH9JgVcbh
5psp/AmnEq+a1xJasps1kD52EtDZIo9gtQ8H+mEbg/pvNjVMqt9taQjpxngPjUQewWEbaC6LM9kD
CeBHenicruVoSAFNY1uWDsp5CBEjqGHtTSkpzi1HZ8aR+hwBhynmjXlwKl8FS6Ghf2hdFmYcCdeC
WpT/X3a1R5zC1GgHMGTXtyEkXyal5ZoYOs70TUL19zhYlaL7lzOrLU+nMP1xKYA7M63K6K4miQHN
9bWe8CmBX1dCnhjkZs0VS75DGsbv5tLX5OMaR14c5mhmY4Htp40E9IsHFiCE8xarl7UBMwJ26FgA
hiRrX4qbAKSk54TSXvvI7BOIWdPErNgjNuuULpDDCApMC5OcNQi2g+NhBVq+O4cBRCB9L+YMT70J
sXEU0OP1hkhjssCR7aW0JPmi5oH2R5NQXCKShy0sCkPLlAra1fvXAhHU9vBoj263NLb5tlSDQWza
DWJUfJ3WjnaGRUaKxFhpqEnFCTL2tSi4NS4yO4SKi2hhiuL1Ozp71BOhGPxci+GEIAH4jUhUQOhl
1l8+byLOcvglCtMLNDhCxG6CQSTt7rZ/yRA3b3HyH9kt4YTKboINm2oqyz5buew6cgJyvPJt4BfC
SHN/pq/VYgdj5n8XpX70+7Fau+E+z8Mr0G+Fyd4K/8bLYEkm3CA4EY9oB0pSsR4n+FQuSMjRUeCT
NTMQQpfpcwzDa1ZS9a9mFOEu3n+fJkze9GRPAUCxMj2EKIil5f115TtnATvBBdujKC6t8AJLdL/l
jNH2gfdiSLtHB1QqltRX1Hh3eclcMXanaRnB0H0vTWsIWtybXXHz51Df0mRlSlJXFNYjfMjiq5pd
qB7v7+sr/oIcEYE5575cMZUbEIrnLkwWjgUhGlBbG3zwBU0VHz5UgYpj75rVipOStUf+3rxod8Z0
vql+EOceZ6vQqjZCt9JWckCIbZZqO1yvEqNZfvTGSPSTw3+N4xOar8+v7qUJ4tDxQBXlHF8B5+LI
tBS2WGSQm7S2UaZaPkJ3ORqzhxflHISfDYXbFwPE5T0dJoavNeZKK+t+QULJbRu9AbZR5QFvoeqZ
//PgxrE+U2UCCKvTQpKuW3hwfShyIFOInJnkFZ3JbEHCXEwFRktz21l9HnsxnEfxPadSHq9+I5g1
yMfpEYiiUvuItxsXB33bDoncMZvor674q54Ospr5ctvWcNdCtR/QR0fLQODLjX3oKrxcPqjkKPDW
6wX0Z4PCAY18uhGSRzhIGqEn7nkDhU0EQgJACEZj4emVlor5eQRY8YeAn8p0MPwx10wBtUtlL+TF
/Ib3ImSxaTXnlmKnwklX9HVdtlImes0ucpp04LTECdM4BoOP20FO9ofLiLBzN/XocCSYbn/OzFE0
QrlPg6BeH0QQF9kptkgkv7LMirgp2uOlMzRiQvVrn7uqtTCogDcnoSnWVCwdheetDM+Nz7o8OOpl
kxLcAVrIf/0YCGXlksze98OF5C9Wpk6DvFV9Adp5VNapKBAZKD76/Sk9/kS828LbjwkEnCrh3HWl
F7LRDURQymawwNJPHR0kQyqqS2k6Q5N5dJr0h+nOdXHgOTFLBsVHGSxRvHlN/lFnkbDU84fEKkcW
YQVIOVf3d4fbMGAOXUEpRRVav2tVbWfjw7lujcIH20Auf322EvK5sUrCexRhlg+3oIhngMlO6Ocx
BmKbp1/Ja3nT4lsxB589Ve2lRKncrQP3Zwg9kBlYG9xQ1yzOPQ1E1zw+4ph1drClf9XyzsUD1HcQ
54+LR+aK3+a4v7RDwWE5Jg43LpLJ7NGToppzHWLFm/dx3vozNHQvvd1msM7nWQ7y3KaWFWIXbkx4
pj9A3qblJr+vBJYUUmJZhZpGXbHHdvhsKoWgTGHWWidltR2wm5ZneUCOkMoLngmBCzD0UgBUeKIS
yTYzoWdLVZdeCLqjx8WejiNvpJTv6fjWMdjNapygDDHrc4zJx2ySwszuaQDf25n9ZupT8Cc2V9Un
2uwYkmvJsL6hkxKds16iC9rDABrQyNF4SSLTSKRtzGBBbdogBT2X8gEeGtOVmBLoGxNOMYdznlw+
grxXCEW4yLReFY9WJ53068A/6VWgqZ2nkqamsadtgf2Xiz4KVabKu+Trr3rs8mIqP8WjteycOhlp
WaOLtNAvmA4wu7z8j4QUJ+ZxcpSnRQx59qGEHqHRUYzxzpLyO6G+zG6aW+mX4WlH6AFJjQn0ETe3
q1dnpMmEzdiNoTYrCxCH4+bS0C6v+kwTlhwHoVj9+GLQsISUSaWSHG3CHsOh4YekTVOTBwPWY3eK
likuKbmdx+EN2ZamOoYYXO56sZh3Tpky++aiUWBZ1oHeuv+dIlsLfy3CEL9Nx1xCJBcce56e3RvF
OPrgmVsw4gbWWGTrsmfz78cbrQII6kRyzLIt0fvmNdpJtUxAauIZqiENuCceuBPr11LPkOPPPYa6
N1JxvnJjgH9r4fI5ANGafs2wkBieTpcCljhORRyUBwL+14P3ekMRSK0WFkDm3UIvsIdowxsxNGS7
ubCw+M36wSn8Dh8osZIq+ihwGde7YbDcextAlzQ3lyPjU9uMn27kPXdRBa9tWGEDKScjB+Jtw7IZ
TDIP3ZN7NlZIjnMq3zx54uVM/CVm1XaI/HOTiIbUF2oL5KBp/otN0G3bFlQME5iQ69FZsxypU9gz
g6dH65VU0rtAmGNxC+f9cJEcNGlyn5yf9avjyaZRthqdNKrfLaYdJHGCU6GLr3EnJ/tKRsaDY8Rh
lHe8DdFktZORS23lPUwvWnl0j649YSZxVEY/LwfD5YCt6jVP3L9vclt+Z5cRnZkQJMk/S6CQ7PKO
LV53qefBpSDYdsIzmpMnh6HNObj+HNsPpTEIuV8mVW5OPKorCN6xP8voiD9zHJty54KRbvUnZbfg
H8xh03w8EEh3d8E0Nr1UKgVJzZXG3Ys9OTYOlznCUZMXYTCIw+svjVQqcW51nIGdPFcjRbp5sR17
+hMaUZnGIxzfUEeR0MiUBY/NeXOCcyYpUyj8qxkHBZlqDarbd2u02NeDKNVy45suipklWB7gygu3
0mhfY4mU0TWou6YaxQPtluCMzPXYCRm5tOFriP2XJsnIVj8v1sKTPm/eH/UdfuOow2E40g3EocVg
UL/H4oPGYGC75wqp5E3hR1taK7iGqBkTkMXZiFLltczTPDQHvx0Ng2qhM0ZKNH1syeB3AX0/7Lxa
DUGqOxje8PJnW4wzJhEVmFLRVY6V/BXto1LaAx2gvGtrDds8/HzRR88h2G0ZockpaOtRodsZhDWo
/apnZ6bNbvUbm5p4ZaY7VIPLCbh/lieGOL7WTEdmM4B3cg+54UCni61NoyY4UjhDte3GffclpYb/
TQWI9vqPiejrtfmwVh1VVYS1xl8QvhPdRLCPwQXkwQJt5ZszB4/Wxk4vdRwPpojNlmwqpXJ3289a
C+1ZcdI6L8NtE2TobE0X5l9v9uceuiXyhzalCTm7rSaXKR+ZzXjxYX+ugMFwMicAZG1/Aax4aarv
Li2PNci2vJeNJMH9tr7si60T23zcRfY0iU5UunlnYLZxnHr1QDAhrL97hRn2OGbGlMADP9G1Hj/V
2gB3GFeQ4Simu9W0JSoenyoR7T5sMU+3WS8I1neGhFqaCeQkiJwrNwox8hkl7mw3mlpi5RLelxS0
xUxSPva8hT+BT1Hcsnux0+FwO//FvpujBdBnba9Sd5f/J9hhWpNNiEd0l6ZEZNBoY+iNbDMS8d8B
CZNDBKsRt3pJgL1ibHS+kPUmn5AAY5kCJ/Vy35+j+Kvq745Mmhy2YspDiiy99Rpqa/AtSZSlkX1g
WBJh86Kg95MIllBgZUmi+spVlvj1iCRWzfYMk+IbsJYwOi8VrEFjDiXmox0HX8dvWVd8seBidlno
uki2sGGDPOL7Vc2dhTDzAR1Yvp8EOkoIlDHDbsbhb89LlGrrCmOlWa0lT6PqtNfN86+VpcTuNxAh
ZqCt+H12n0KNzko5Y/jkoWI0OXT7048XDwHC+fZh05bkAZWnl26WakYaXeGbSG+ABFTccFv4anz2
kI4kbEfv/eq74hjG56rFpNhEAgESzFz47ezFg0htZrkJXlj9Ym3MMoHWYGiaRQxanXR0YLjZwbzY
CIljdKYk/RGCkjUtKxngRlYfS0xHpRbqr5vru0gKk3zwHMsAjGIchAQdF4FK1qSWpdvhRNYhD3x+
OD+BDvIZ/TNIcmHPcqOoNFbXOIL7/k8ypd8K0EjyUBDyPq93gmFbPoHAl2cPHf7tPd3mS4j+iYz3
pmTHd5Yi2NLS6oVTnmNvPLe411Xh3CfW12OXGMheqv7+9E5P2wKu6LoGVtcwGRZPpyt3hCcUuXbU
NlYcpTZWLfSyRV+MQbNHMzf5dPJDDxWUUFwpj9oAfUCZ9PVCBF2RR6tUWamjJaVluh2QPhHDCVnn
9uGU0bh+KqyU+N2C1ItM7wd2xKQj8fYEX3qxpETiQNGYfqBLFoOGpvzihIWqiqWFETpqXoZJDUzi
tKzGRv/LK1k09TJFJHVCTKeEUv1TeyuS3N/FrKUgteP17S2mvgx3LsPlraF8EG8ShySWPqsk7IY6
y2TVpjSyFxC16vy3vMYCfRxebjbNPnqNQ9IrWT7R2n/uik0eEhod+7iW4I/F33Qjlabtl2x8lz2t
2YD+J879jsPnmbI2nuCQFy8XIMVTZHU8frxockdm8NVs+FxqxfKQhKaWuby8CxwOyLmLd2imLpma
BGom+vV3ILKgZ0zODmQtYw9MWodMGL/CMi91L0AT+YD6JLg5KxGXAp17IdgkimrLcHLG6j0/Zt/b
xiaXcGlKM55HemQE0FPOIH+9fXhqyToRz/OanuRhqURbSiTBEy8rmwP08obHrYQS/Oadu5H98XTx
FSAYeDTEhRoP3gZVNfnuvu1QFNa6s2jLOpr7SG8/lfvhWHaVUC26YKJNYu3hhzIy+3Zawjrz9tQ8
Ylqu7wtddX0wc7/SnJX1iG2UvWooGIB7ku4RK/ZZAR08/gtnsX2WnX9kc5yeXUb4FdmDFXhzU1IC
naNBTvFUqLdFA1S5MvkwDX4uon0ZbmnIQz3gKiC53/2gUwca9tQMjTJoqxJWMPN/mdD2hKjtgFiR
RGjDZWwAk/uqbso+tl0bloDhF7HkaGZ6j9nr51tbR0FEwSoSwiy2XdtBAuiX53jJwyqZ6HWc7L1l
lyGfUfENk9AVP2FKG/23yCb+WkYeDs0MufwlLAOsGo09/PNIMpHEUKvjtqpSZcYZq41omR5sJXHn
hhQNa8jQw7C9MuzyfQcJiAoIQbr/Tp1lq0GGMMpAa3cQWRSvfkudaZ8HPhqdXp3nrKEgOs0RM6iE
k7h/j3dOS0bLfUVM7+BBdecQMX4Nv8YMte+2aj+1DNpa2ZkqhWnfrCmm4kwRAvG0UMDMze4sSqMj
8A9HP7W/7ARAz/0mG6FyK2nHgIJWtVXgim5WJypFvWe+bR6OOsJJSN1qGoO/Ydi4BWQCJ8mTUwjY
4JkkqN+Kf56FeyLwwzhnTk0SDNU6g1rqaT51yzrevHWKCmpHfhqDX406QdAi0sjpU0HJCw17STWL
7jgLsDNGLvTI1Em1Uk85TThmMocD3OPy0fvjCxzLgd2REzw8dNJlOLpCSPM8DpkA8zvY8hTT8Efx
+FOfH9duGZdZnX9c080xpS8OIGCis2kYfE7pvAkNV/zljGmrL4k7lrrFTC9vpvMUAc0AU0sL/G2s
BQ+FdgIoj/rWv5ng321eNmijHdkxsUB4U85eA24pTGxLotxWGpEbuX8h0H1c9dWtkJxKGEeMkSq8
ppFAcUU7zCc1rvkFMr+incoP6Uo6uhz7CLJ90R1mXZXjHYdF0afZiwpqJIyq5t5dx5Wg+LwaEiZQ
9TED/+tyOLtrfpAmIXM0h2VwXs1Rq7/GxkMPzAcgCTFwWR7PcesicMfOtRFeawQ44ty6SHo14NSY
jbXEQfNd/XNCvhXsIYLoPNAB0wRkndxOSnL1R7x/CRYTqbWUOMtcbhKCJThxzq4U67BbIPI1WWCr
A49cUWGQJj1ZKbYRf5P6y0+ub8ckrhor3Hpf8zPRZ0PaZ6d4MYbi1cRkLaGyiOclX9ump2DxgH0c
QWDl6NCJ28pAhLyB/4GQYrTUgORvAKN0lcz7Fb7xzTYVs9YkvZTPC03DTyhhAlmdBvPW4vzrtIGY
PLW0/RsH4lA0bk/yptlH+YFkBMjIYY6CGHtxOV1wFTgg2skb35RC1mABvYgy1EiX/xiovLmSrJiy
8JALzALvrpqxD/3eU3Rutk9jLt6z115zQ5xh5xt0GtsdJQQ6+wWS4MENOrPhyXWv08as5ZfVnE9Z
OyaWIG28f7FTG0tKe/F2JdyIc2RctfH12k7GrtjDwxI/SfeF3jScIJKktRSIZlFAFmMLMriIwFks
4dOp+LTA6c2mOeZpFISL8Q//aDvNOBa1yijMBRGx9K1cSyrZT1uGZXl5iNSuq4qoHByw1658tuhm
F6rMonKG6SyYG5lTaAyVVVkfmsRcNYkyNt/8YePi+YaanshJsb6/ktZ6Dgk2v8siJ0I8rgxhUf5p
j1y1af9kIw7a/9CT+QU2NElPwo4T47FYsoPAkOt6MUNR/GJRhbHWJmIoMTXxef10qt0yU94czbaE
PcpIfOAJETxoIp6FGaia2/oNlQHcjZJ8g+V5SQe1xQ/mYpl5Wvjq+LoHa33GRR2NkvTfBmknckrd
tEIBclPA0fuyyJQhGmWywZBuGMPsjm4ZwcMRmUL+CEZ9uA1bEiCGbPUgEVkpUOOtkcD9pZUo/93b
83YtBgn2ogaSIAJw+8R4ix8vnNEo2amdfW6BoJOy748vPtzNgu7ZDNi+ddC06gILbaHVNEfyz46f
9a5vO5OCICMdmPCAUuxSyaiHMzt0p5rBxtKfqP6mA7xK/VIB/8XNldT34TJq3ixTz368+GNoEwZm
f+hnYAVU5GBu9L11NG4zcNGkcrSO9Is+J/NeWqvBgm3/lrmKkPpL9qCZPBRDxywsWg2oFAcj5+RW
ITd4ptMjPUBzj9QkcJMzzgg58EtPKnJplcuJlmOdr+pliQ8iT5/Ln4pdzKmVYemhlAYWhITBWaNC
Qr7yqlrkpgxl67gl3CCLfUiAi3Wteza+Qd6yCZx+DeJYMtr8xMG2kBZyTC7kv5gqvNfdTHmSxe1p
gdn6i2BEA8rn5viDpJhPM2WusgOachDzVoxgD3vj/5hzal569cSE68cJSK30PQehsvkvlnwZ6HT9
/yWwF0qrXWNNvVvsHR8Wm3URF7p2TjlYcmAfNLn0YZkM1ewMfKyCai3tlq08aUs22qTQDF9UUO3F
AbM2weAMX2MkJH6TXCQCSAcjhdNG44wcBXnUDTQZUojc9blhlRaW4KDiEnC9HHeuMKP6Z0Ku0YfH
k/NKZ45ocWK4zIlwKgckwp32SKkvMhFYmFRXJvXZkUivEGhRgLw2EzRIAOp/D5nigmH/rbTIbYf8
v0r5cuE3rMPDG64yixeKy2bp868WHVHrKeb3icK78sr/vyFmYQHSAr053Htt/1K28GPUUIzAtXUG
8ILzC4PFGrMKuBO6herXHh/VIgttUuCDYsXTZEptL/luNxgaB1tGtdV3IVpTxiBLTryinKZSkqpW
9h4QOuSNjdSGGAAfaxYMHe1eU86lCeMV3rZlypiU6TxxdT8H99C7CHjmdhya9EnrHBhMi8w6BoFT
EGFrmhwj3czi+ZuPWKqvO9mC1rndrM+5bS8uumxu82/i7YfFRqpKLDY0SDU1JXCu5SrKda3ljn4n
7Z0dclHuUwD4t/AU1iNwvBXUIUBXQEVE5uukD71wMX9uQiT2uxqFJVxKw7vWf+iFycjkLXR1ecpN
TD3715V9f/49uEd3k8a5+E7hWEOh/3FaZgmvWvcOIQQ1Tsl3haRs7ZG8luXoa8SYdtpOC7DajAtj
GsVNVl6/zA61YAkQWtzJQRtbbG4XCxYZyky2PqUiDk39JBKaskrgqSwyaBcxYIk6b76rV+Z+/0fb
CbrsAJNHFcc6yMn0aOp4webX3AV67bXe1ICqx5B8GNEtbZ4gfSKYk0a6mjvPxhfUJ4h1wisJdaGR
gjKfJYvB4iMA72ZlgZPJXGdh2MYz4j6QgKQBiLhv7Px6Y1WBny0EI4RPGN3UxAws+VwIK9vOMqz1
GBTP1hp4Lvj38nqxJBm0/VcWolMrAa8zUoIogHTLd+5IalpbWAjTMZvFcsPLz9Dd4Kfqe7mRlW1/
IXfcYW5nRNE3oICW+rY5urht+q7tXE3gZ3CGNFbzglX9Lw7jbrHinrGF0yHQT6qXEtpkIiHwO0/s
W/YWoZiN4gTuk+BDkue35NMl7qunR1+4htkFwybgom88olL6x6vskY6z5S5ALkfYpjjFy+Mc4txt
SAD/dmzXJojRqKzL0TaKZFP3yxdA1vutRuoxGpbqCWfpj3+bKMp3PL1sSo0NFXNap4tki7pd2/pe
DZ0m6YwMwwfaBkFl8vWN3KHycQG8epVYDIa+p3EsraPwIrmjk3xVLPjJa+GVqzq+iGc+f0ZVZCSX
XlvhhYYFSD5y7jZTBou8Rhjj8e5HUjGObdOKGL3nx07Sz2E72mzo0H7dV4b2bXnYi52GlVBR5hK5
65GzxPjH8KgS9wBf5atbJyRNb2DncnVmO7cpYla485ZvvAnxXM7rO3WSeeLgywT6wXgOdVeS2Wef
3fBfeyR5lZa5WFEhdZ0MJeyWdMBeeNdfgn4NvWh8HzlxEsqfI6+ni3NjqWV7AFUjtTMTEe35QUHn
U1viux5c6zepoDXfAUiNuMDrIwe/W3hKFSCrrsyRG1mHVkyqukRt6KxBuQHf2nkI5dT6O0iQUabZ
rvHhaTTKwsaEJKX0JduyZ/qkVFtIktFDlAw2c4nVmZvuKsgu+7ihS0xefVz1t+0riWjCPyZDu/e5
/CcKHNDiwSIM5/NY4tPXPv+WeMvynzbxHIaL2eQbbkLTd3W7Uz9qu5rr+C8ykgY07A+YPRKI7fwr
nF50gEZNji1hQkcN9RKQomKmh/TwKEvfpyNsUhktULE75nECYYrsHxwV5jjKGjdArPUvoN8gbiwu
Ho9CLO4URDGqO2abB5O1UEMu4T2fzD30aI8Ns5dLvnwFIVjzkgPGpBYfEeCPiXtZbMyRxi9rU6u0
QHTGMiUHglw6dLuvJTUm+1bbf+NOhxk9YRheiFcXvcgJXo2MmZkJv5aLe+2y/1kRVjAhkSbvVdG2
mB5g/D4qakX30HzzW9AOs+bg+6fthQx5OrhSJ6rGlTL2RWGRnNsHJv8EqSGpn1acCu17oQ7iXbw4
jir+0AE+ErbFrLc0aL7auMn/gl8X7leY8BMLpt2Yh/WgMipF/CJsYVPYN1LnHDFEmTBBgoq7Wuds
LesQxeFIg0dSVNICHN4L44J6dcI/0W378Vq1uKSGA8/IEwxIamc7iO1gRhi1HRQc7YFQyptSli+h
cw0PBwqc24R+LfzLlnd8drQV2PQ4dEj21pGiX/7OXlpFsDREOKWnPiikN2kMbnmZszU90NfclASw
761sGawDyFjtRO2qcrNX0UbBNs9yMRzk3aLQtQw/JOAl48dHIwepQ1dbxiZJkdMVEqWz8U7JGJAJ
Oz3a8YY9wcEwZCZZ2KjR0GF3fk/+f1eJuOK99QKMtvqETn3RtRatSoZm/aBA0on2fPE6MMqFYTQl
FeeHZuQIbrKv6iTHCEjDBDz2AGZ4UTgu93mkl6IiWGHUtz7jRWg1+B4rkWzDw1rkMMpyAX345XB4
lP7ep8IJlRTzTRYwahDps4wd9W0vIGxYaKUek9qdbvKSLlGTRcNVU2FZ1kkI14UCtBH7UMM14DoI
2RHuhf4VC036qxPCIAq6nJeEKdlLoERHP0KBvCLlClvuVNtCbcp/4YArn3b2wK2G/oBKqhN49E9J
silUv3mHtkBZX66J7uyy1KtNHFwFlXyn9e95lPyCAVgieoeRrg8V3lEnkzHgSLGIO6LT9oZh7hz0
SaUkxYVIqKoUITgM/Qp8FDYKqMCdaIR906KnstKdT6O1SlwY2rnwo1ApQtB1yRXFzolNeUrYdfjE
658/lrVA0gU97DNKNZgUMPd4iJlSpgG+3rLZHdQfgpY6V5ejMs0LfOZZU9T044XY6LZXoZmlbJue
IygnJs2r6Clj24FzLPYoC9U0eO2C8UjuIV+FvEEvfNgSr9rp4T05LP9WgwRntcwPtRCXInrAsL7+
Xu8BGnvr7DCKXiZtpsd/RzCWLFu4CG0Xrli1PgSLtQmlMWR6vdn4LqZtcsp7SZbnWF9KHvAhfSA2
x8dTqBd90oJTtEnbjEVaF6JICfD/iNmv4oLuPZDYmqvAbpIUh1FEUXzoZptNarZIYIf0gq75tLwH
VPhBQ0RAZZunPVmblI/F/0/0GIOcxFsAdcPhYHbQp75w9AGGJTkDwWv8rJdurjVdGMBmcsKwmsrV
yo8kGPohwayRXTbfgWLn2qqVxrTKSTQr4QLD0rLT8w62W4Ya+bjQDssLVk/ibKtIpMUEviL1e3vu
BTJ6WyoH47AjHOB7Co8jz7aIck/5oxRi2Fg5sxO9lpmqECsipMS9PDJUvGLbl7JQX/BJbZRw3FyI
wc8tcYDAc6rmjvWiE7bOXDJBxIL5CZftHGXVuSQzMq9I+Ecl0MeCGTZMq9HZ9qJEGWbVsPxDGntg
11O5GaQtfWZu4whu4JxVh6TrM3xARDNQ1ZfUdqhUgbu+hXJsT8iYEGE98aopxtE0iscUuYbNTE/Z
ly6k1vtNtOhq327wkHvAQb8BA7cYEZxIca1WSyZe0uxT/J5/uBLqLoUXXUzyEHC+FYzpWqcOwYZg
IweiAgZ6Zu7wFoPqev3nXN2l31xIbjWTp7l5RxQ5rQaUV+Wp0DBgnnQ6vxsvryvul77BwL6MFWHQ
5iBH2cjPpNVysntlWlvNsFhAS/YNLU3IJKVPU4SKDWSl1e4pCEGaA+pr2IXBGjzn90KLx9529Pu2
vdpZLhVrsEYeMPUdFqfY61pHJ/6no2rGc9NcUCqN7GtH2oKuZ5LHUxlIzkzX6E/S1MghwYH39On1
BiQzJyuXgJWICnQxNo78qEfDLkeIUpyWZ0ZfPyTb0AEHUis0OosUvCAL8/t39VAOG3pUVVl9DYgO
wgewN7TehmSodXREvyamu1oT9v7hp8twAV6qC4/OkPZOG+UeWPMpP8q8AJ/Vn+QMqHhDCzql3wZk
vb0/UgACc7G9ctRyMCrlP65OXzQ7EvDcVwwoJCtBNOdGf6OcCiqTxe/tx4BoWzC5ggKuuAg1P7tn
fBJnNPEI38JiEKaoDDV9bRn3a/Si310oVtOGEEqkNJwswl5LpytQtUXbyuHG9GyU6AQNjMBiu+As
En9w0Nb/568lXK75/EVup/N4s1hNGlvvPI55iuYZsTAIGyWfvazUBXyd24YqefWWsZcYzcx1wVOe
MUh6r2M5sSDi0DL+PiFVXW2c3o8haDF50JIWpQzjkHwSJC7+bYPKb/79VhhUfVz5xNx7//SGXVvS
xeTAKwD4NrzD3GwZ0kn62gEEzb6N1QD1/uB/tX10tu5DFGmJGyZ55z9Rh7OzgSV8gnhgM/12LrZu
vJXYvTGzlBJsaB0v56uWNUCHRwkxrIy0UnYX8t8G8UEtHrtRcb5b7f5jt+7Q1xgnbQ3nQMNG28pA
us4XNdTq22+uJPRjGPXO9+GhGhM2bhIMlZGZ1brQFy7JObk4Y7NeepxazfPcrcP2G90ghKhcck4K
ZFw5IhLVFT3y1nbyEVJg8qOPYUYBzNuQjyxaOvG61Htiy5E2KupX5BrDIKToUNqCSRFLVocRBM0y
sEluUX4SQBsvbCGaNBTPbZi6kMGm0GGh4BuHF7UPLpASDM0Sr+GpzJ/AqAm86yk8AXxO0dQ6V+es
LNC+FWG9YJv6glXH2vbQUNXbjJg16xFg+5oDG8X5SkRC2oEpTPa4O6OvCZ1PZ5MLQujiNadb81X+
9u/vm4EqSW+ebS6/9U4jublK5mMiU0rL0EPuPSQ/5Q3HkDprpQgYHae87LP5+5cR02QyCHuaW3iC
RtJYvdn7JLtkdcjJycrNVqBCckVK78vBivo1NQLeAiDsHmg8VMPKrQxDgycCUxumvjO7AmNzL2jF
yKsvgrAXhoDqVIVDb+PRbHDLBtD4wqNfHWJMcHaZmVQ2XEe+6M94MMIycZ2NN1joH7Co81nWm1pv
22/KdbSBDKSdIxnMKQ2I9QiE1aafwln9DLzFwuc+haC0VOOT7wvNmrx+QD61iP47rdkvzl6ZrMQo
UTiec3pWWl7fnRDZP521pBQbrOShaNEBFgfVqVFSpJIxomd7lipOFa+RSfRp7FCevStkWfMhrXw+
AU/dc3EI4OEW1kRyfYO+nOBbGJzaVUMl7lJawnPQfhicXlzDQ/RY/oKYuLHYHanGBpKuhWY1N8W9
6pUL98z4GUE8TRwjHO6MHr8w7Fq9XsScpT5wt2xeYQf3A0bf63MPmnvA/rdvKI8cfGlhe9JMoxH3
3h6eLzTMa++hNSiBzsfK81D8hk6jFG+3YcKKaiInvWYca1c5Lc2YRkfXKSTxFf8LO546dyNeR9cZ
AFTi+3vgsngR0zEG9smlwx7TmeC6avSeNPaMLN9odmdFeAQ3DYTajozUNiHhlVmTsqpxTcdiSkFZ
uTCMw92B7EI2sdWD28B6B924+0lixeabSDp7l8nFNLl/3YhXURIBz3qMi5+fRNChXFoQcovgcs8L
aS45PyfE+eHRn833YYVXDW5hPvbHxgNUrAXYssMG3Eulf2LS/X76Y4oc8sdHjBtGghMdudADVBw7
J6PY+NLaOGjrVDP5KGoJYPu7xOPBzxZ8ZSJ6/XUX1A2VM7BU7hGbQHbz6D1s158gVO/6/0xWr3nh
R52i/je71632UX4IK7PmbLtPmMt4pTfzdtzrS/OkcOpd/M7hCkfvBrgaqIjv6U69SVPIBsRLDoJF
c+faky4VBBQj5NxWeH4r+rrnjgl9+uofbt24KXgDJxdReHh+b7aKrUVFZRN6eUAQ++4c2/NmCV/V
S/+bk5A5oM68KuMtaR+sG+iX3ATuQ2Zh8rDx0rNH9ZRzNz38GybBG1CMkUgeAlA6u8Qm4lHV47mB
ahm90HeDLaOMpQSjEfBVapGotrOSrKse2PiJDYST9DDGb+6dQnv/L5J9WA8ALAOhW+iWfgkdy6zP
sFBKqCUy/mO3WXTggQFINP+h1ngkwt/iR+lQaeJWZGRZ1npKLWtScicixTlWs7CaESr3eURCk8/L
O9I4/t0Eu6Jw2Wm6dnXLw7+peiBUsCr8KEaT6bfrY1k/bBsISVMuwCcYuIaofeu2m++nFlQrJqKe
H4F8GvG2fv43X7dVBo1hmHPDxFO95NYfZ5yINIkWVeJkq0iDSJkLAWOVu+T3hJB463SUUD76iMQW
OIgcG1dapwYNXXyK3gYXeVXle9z+Sd/SWS5H3uFcQvxP9UE9mJMy+RmgZcRYBBkNMziAMkL5YHEZ
Npql4ZLVsS9eRTrGRpIiZQ9S7YNtjDU5x3jCSQie3CTZTkctmFiNGPCcxpTRAjUqB4pCFytWTJGG
wxf7mZrpVzUnsgWonBNlWakpiRW05ivLm8VMS3Bl7H+Ez20KlJ0+xeh43IWTBCZNyVhpE9MmIQag
wP9nBkob2MxQsFFmNk53mdl/OpFBM1jm31NHvDAVI+0P5PLk3ZxJWbjt0xeSHmtf6fAK0PMe8w3l
Vcj0353eEEMnquOgDzfpD/8W+XC0fFkaHCfs4gWmdUuuo4FCa5gT/Il5KwqojArTP2nOpxAwHbdm
0t1ufwMWLAhJkI2R1uE21q13YOqKYzbwGzzvf7/V202m+UO9JZVB6BmmqJpxuDFj1IU8T+QWiyqP
UiLPO4BgYs1ngiwGoaYW32IFnG7L1sK2TLqxOSWbJRdCFdER5/jrkbIrWK1OEE2ZA3FVlTnCn4aA
1iV/HjjL9yeZ2YsLU5+o9WjYG8g5HwIva5Flna8Eb7sDbVJs9klqMDPMt2kca4zE7CQsot1ojHxK
i9Wvc4Vb92DvmodPT2ytMW/W7hgq2Ek0iRLdV201O5IQtZWiIVxw7fQ6c2VQ4Nj4B5CSo+OWjpyX
hR9nYJ66rvdyfMaCpx+tqB2uveQhOrEuhrayhSR0uFtN0zfJsS1JAIMuCUSUvkQ/QOuZChADtL8m
MRItSqFzKAt2qw2DlXeaVp+ghcp5bcRm2cFMzrslogGztwq1suu1pqCHsYok+hx140C5ca3hPg0m
SoqnN4sNaLzwDK1Af3HzoyJeZa8C9mcjPdgrDhh2pDSEV8aPW65gxIvc26u3IyHu1HPfBsz8sIN9
lvNrdoK5qta/wWD89AMMu/F95OfltVbCtsKxUX3boln9CVXIT16sxYeXW17VqMzy6mm4TM+TBeGX
SBG2Qt6WWZfw2J2r+dv87g7jrBNnsrNw76Yub4E7MzoPl5IAqWtZd/rCXXWXMoRYIQRRLKDvoEDh
mWOcdLyj4RRN19BzJa5VrQCkF30RoKq+KGONqechRalCws9m+kpXUFIqh6ZGC/IYHSXObD4fUZku
Hh6MQWJn01IoYk8Kii9JBqjen99MCDZoqEqS0ctInqWtzhIEyln/tSWI265US5zNHTIBwQdBt/f1
HRMH6klXRfmqOGYWnj2q41rUaVTfHEMX4QCDhqRYyTdogCTSpLl1n+MDgWtaYmHe7areWn0tnf3y
LHCzQr6WRtj0PBMZTt2lz9Oz+6OlvYyiuKE+af6sSyJ7Mxy1Ja63m+GovUoEJDU/8ieq0wXIx9NP
cTJgBv1APiXiEdiDM2lbZPQl530A9siABaL7tse4yKFVE2KQt1/Esu3HKGonLGy+uA/c8ymkHc6u
Euc6GEZjq12OUp9wYVZpCKEh8bt8mgiHjiTVXJL8jtPAMh+4oC6HlSiF+mjFMN4e2J1iDJCCAx6A
whtv1x/fWWG/sJaBliBVOjixAemSxNL0p15qO/s6/5fxfSKcepkw7UiMekts9m+1sMC3VymeM31C
MIlQkPZgqv4MXS93llQv7m0Mb9Qwc38Tzt3eblufEOdGuCuy+Rs7vRNuHG5kdwxBw8cVFd2lEoiu
k/Er72TFNvLdQ1U3A8lRI4P6U+4jsQojQ8fEnxA4Qu96b7GJOXX7tNDW/pUcowZquX+tmGCpvOM3
TUBO0caqJLk3oo87rMcwu+B1D9fxYVyLcZ2etwiLqnfIsVAeqVhjyIa7grXqAq3nVkndlUVAPA08
wMS1mZzzGJzkOibm27tCkP57wkbTjsnYI9GV5kffwsxwTkofLDxIXo47f67IhIP9oNTmEFn0nbFb
pbl509s5ESqiTCzVE/uPCwZBSf25v+d8xejRhlC103XeIwDB6cazhKgC0ryTYyi3lPm+/bvRfLkS
S3EHpULzH0s9HHZ7QrrVihZN5irCMvNmBoFeFFBxtbMA+FSDGaFtfeqD2MpOeaIsmLmzKe9zGAUu
mT7wIOnf5mbMMJ9rCM0t4GVoDjDu1ondql7i7VL4s8bGKhd70mrvSEsk8wGP2Ga0q3rtoXdBJty5
vWuJZEpmCHoU0LcTLJZK9qie2wXFndYch0ZbQgvtxyF7IcVGQJp8dtVtsV/JM+fslzaKVbQfjbhj
L1BJw4t10rHKI4dn2PqXu1dVkLG+liOvvVP1WSvRltPGU6yxfQAA9xYNRAu96klVxpchMOiA1VYG
U9rcLLGumXwexkUaQKJahXY/psh7ZUCDuTcTRzJ4eFoSSzxWFJ8dvh1bHR94S4uNrKUwlv1piDfR
KcxqSgB4b8o9HE2rOkCjpSrfgfHFCTHR7doqTMY2+uGvcxb2Gm6IY0V+Zai6Npa7xG6vNCMoA/46
J+Vstu268ijFOkgKdp1Z572ZzO/vcHw9KuK54NngJbz0TT85YWqC5bFR5SzucJdsTsCuv4/zsUfo
fVBxsfuJ9u0s+fj4lmgf/lq8lm49UYjfsroqBnk3Kw8wLHQ6LH7JCa6/QuuKjGc6WLoR9LpxvOpA
xy5dFE+Gxn5dbxDScruJUe/ryRTez5W6iiVX8nbKzLlndPU8v6cabDn1gmr6FITtDH93rwUT7pH8
J727BmF7WsuXs42F5396Y58FwN9z3VgiiiMjr6sNZF7oqNitnwzcZcknCqc1IvrRZISntrlCkI1H
aJJPbpD8sWZZ1Qy4VIihFlIDiQqMf/OIuS184PtomoJdwGqhDhRCxw2rvxtEunUeWuhAL/7x58Ql
JNL0ObRx9esEkrC8aqfo8MsYC9NyT21yY8FqzdvdPSYOXleWKkeuMRnya5+embxzurpPseemVlAl
fNNtyEg+bs7TXH8xh6r4806nZ6aZnGTuOr6FaDlIybWzb2F8y8zfanokMIbuiX99EMmCt9ElMlEu
OSgiLHpWJjh2DjXcjeofq43DUJIcAR3jo4H5dWqc0yCcfQOaRmpHKXiAEIPR+oU+3h/hWS6BUngd
6UrJXKyLIK335AXxxt71ODEpk1LnNQ3+nQ4VYgFyMF8JAMT1mS9w9UE2SHS+T0UmTYuFNe+QISjq
HRHFmVmMYeBoXm8drg9Zx01JcQUVxXp9ALZKsjTKJQctRw0vw+YzIoEWX5n6UKyl8hYAU/QgD92O
hHRqdfwi5dxfybgpYLZ+RkIV+mQkfTBKLwdvkoMTxZ7zMQNcSZili6A8HogzaR2HJI1n5h9/NxK0
dLeRA+4ubkUSR+2WkXwB9TuIkN3BIJrSjRytGAf7PCiPEkZHqtSu26Ebb+YnSlffoqA6nO9pliP5
HOXH7V3j/7IeHI796rJRUcnpMrLBbx2z4ss0z2r5eFvac+BeQ0KUX4Bs+a4pjm2v+Zlp83xaQCBF
wKz9l8lyNcdxUB2xBvNjcqASLvKyPsxfP7tOlJGIuN8t7B4A4ud4nwOxRDCLjEr4aWsAziG8w9cZ
PJ6Pu42UETLQN1BGU9Hrc62pYzmtTQH4VRf2flgUh20s7yYyrOGYSTso9C5cSI060R32xHCeWFIO
4QV70i/zZS1iB6LXJIJWq53bOc9ie6kQ7eh5ScpDBQ1zsW6b2Vh+nHh0j40Nr4AfjuCPtl3DMDrq
RSWjzTmlPhlE+sxflbXonTzan2fMdiwWmWLge4W2GmOPkNCmc3rOMEQAfMl/dnOiZ8zPeQ3R4e9B
UiNnR/HxsENkbCQVLvU1y5q+jRVz3kAfZmloj3UespiDcIqKxy+k8ul0dIwm2hfhjMidKAJ5ji3j
sAsBtyhZyXmBeRmvldHxWJHaunfP7+S0DVt+Wc3meCx8pbjtWpdJezkOjs0EwBEE14zmEpenmpkn
1Mz+ZLjMwawMApfX05VgmSexvoDJNmtdXQ9t7q7A34kkKKqHNwWRarPCDVRRlBJNIpEa64frjO3M
V2CiMfYRMoNs/JyjKnKd3yy0DnAaCAdBPKnWTT1wVbPRQKJp7NlWYaeIaxQd1GRdst+QKADxXKFM
3elx58G522UjMeqYUvmiUCHJnOKJ+MWI44wnMLkIY9VyIYnbeVXXXucsqBc5/kiRKKAkEkfR8T1D
e/zcNt/SpMDrYqU8jcW0W0KQkQDWMs+bLR2EVZK2GIMznzs/Pt/1SjLS8A+cJm+2Hrn6hnjN5zj1
1J4/I/YJSSXurRMJWyOvokpDWzVTnyqCJgQLGJZl7T1WcT/qMsu5NN9kIiARPv+ZzqmgRlqyiERM
7j0n+MF3K5C9AtzHWUjMzh4yjuOZLmAx4Vra/XsEj2tvROXBCFRDRH/b2CkfxHxauxf8mB/VFX8D
SO67qnIhkjZFTDj2zIPiONT2rmG7qGdI4sxXBD783styHVkIjMaAVA3ESyrnZ7l5sqq9a/qlNO56
wZKLOiUooVTHloXiHc3JZBGMAEcEHoG26zDfQ+szdnvlF1j/YI6rWMUYMU35HslwKqUHE00KwbgT
UXhUboy6fMqibK9S8YRc1RKJUhg7d3UWFLKXWdomlh8i+KbLphRyzO+aa/p2xrEE/cYJimrS/fDP
bcdxmOjIVVRVdGZw15X6T2JoL9CkS3cDED40u0TJ2tdMPQIFcYJL8B11eL6R809loDf/uKT5ivxb
A3bn2WcSoluUNY1VOpX/CW3HWxh6/uOLQlU3gKCjFu53p09YEIzL1CGWiwxdnkMe63dsaQiZ0dFF
9a4zwE06wOR+aBLDKTEY4WrjSFnfg4l7r3Qd0I/3YMvtb1/rPNSnkDta3m4AZIkvpEwlx8HGndYO
P+jXHvdIPl6ObopyA3mHlskMsyfbZejFY+kwm3y5pUmbNsTw+HZIVF7cPlyJ1aPwIJMUP3wxUkos
BhAxz0s/tIjMXEHjjcrDA7KVPWrC6v9kucC/asG4VTsn9zfaHHOMVf7BzK82seobPqSRVaBWEVTu
dSOEQbKq8rrqec2z6oA8/d1wp6b1PZ/f5hT05mc165MdVyLOo64KqFdyMxA/yk8KPoIuu9YQxAeh
dhsxXy1HmXx1ikcIkY8Ey3hgN5mMR8/JbPmZXXs1GveU0Q7TlaHDaMI6RypmQ0MFw8YfCjhZdtew
Wj9xViv88MmsY7zrZcGx+rPKIZXd0/mliwDo1h3L4PZ+bqaWbz9m9shMi8MIo90bIbhWTg2z9jY1
8GOY9topkVtS9BIyFC1jGk8TDAbm6QuvWgCg6IdAnFHEWtzngvHc/qIqBqMT9Vyk3XAHXIVkQWtH
s8gF/oDNejuhOZ03fKIn/ITzVRGU3Kj45zr6hI/lnDmuyZYDnQuQO1rhG9rm6xB/Otm4UG88ArRg
jNngbeLUq423L88bsKRo+KJvJPnBA1O6qbqa6agOYqVFxtnqn8G8xExV4q3uaREAyEATa/llE7Ju
IFYev/+1GRIDtL0WYr+G+EHxsgRMUZOObg2MBowSjRitE37G0kShXn20XFJxuzPJ9bF3vSt6/A9v
0eOfbAWOFKuCu6Qac3JwuyJc//CaME9hzSqLifkesnjVaepmVjX9kMmyJiah0araxxI44AJDGqoe
nYxhVnEWlpxjogZ1G1Mhf/OMDLQ7GxXg+KK1hDa3Fzlx/dEBl+n7CLOWyXKVcszNNCzIWW9Rrmes
glcY8vgCMYR+nnokjiA2IA8GfHJ6gND2EENSTS4+5dNPWbh0RaCJ8bj3b8sZnDKXDv/kDljrFqT+
VinBrRLCZnmeeq0DnbDTCYwer89YS/AFdPrtfvNCe2rTIEAh6QEM7/oYRrZj2vH3449wkqjChUVT
VcqDRsGfa+kuudg1AI5eH6vhm17wW1I82MlQo5kRgW2qhgZB0RGhH9mfLd7nLI5kgNw5cL47zUUW
T0H0kYBmIvqPA4nNhAwYybH1WuRmYKrMh93KsCP7PnpZpaOrsylq/py3kSIXpj8S9Nd6McR9rOL1
tDHP39tBL0iLtURMz7M+V3VG3jgKl5Ww5+6swoiAV4hs0t120Z9OqzJC14oc8MbkstelN0B6+3ng
fkbDuromBh1j9lBZ086rhUpRSgNeOSXBk4/daQVklk4F2B4noryfPERGWlQsPtoBZ0u24eW7XAd2
Sgq9PHbnoZ2keDbR4lxLxtqjngPRym6KeidG6tYtNYEZWQRsKHBOzyX+NtCOAW+LYUdOYg1k/a8h
1b+DPgYpeLat0t4SHUvwdWZnQm1/VLkl40znRXFfVCWfYgmrzkoVXOEqj8fXU0jG1uinhT0eJkbx
Yiu8UsnBa3oLTzvpEEQcrmPqaKoKWdfDWic7xYo10+hscaYUcJVMmzsKoo+OMuRtSGb9k8ehdnl+
uDCrAl39bCb9nv1JkdM+LUjmxRMIiikL2cKtFLNccIZ03uk4KuvHj4azZgrZ3l8p31tXot2rWjq2
3jX430kjE9gvlOZiO2QF4T9AqwtidZVCdvleDpgrbSBocbusOCfgm+LtTBlhH8J45jioOZ/+EqkY
ZkYIUsUxnta0yWDMPTzQRWeNuEGNwJ9kkg3wiBamIBMl0xHZWGAKBuIPVxwMsaFfn+Wq6/UZl3Xb
cskF1i/xHJk5swuY2UEgug2pOLvCJmXnJxHejuGNCMDG4cD2Yl/JEfZj8Gv5xA90VJAzk76u+Xlb
+lpLpmk8C83/RE8QYLrUZYvZaamvSZbU+aINaYz6fTdoP/txjXIKHkfaAdT02WC5DVt0ztigY9Z1
GZSh4WYIJy/BM2asBugBgq3OMm7HRIKXDgjcp0wcifk/504zRZ0xPEm4szniUPLotyNeob7kbAc4
d6B52VioFWPVMC6H3hkEk2RMa60WxlvSTvydaPFkG8z1phQHzunmNfH43cBuahafV4afVopK/akx
bAK3A+1Op/PTtRMos/J4I/ePWkHzFUgtREZ4HbRBCnT1TF5BOywMkmEogxMiEjUGe+IisYD6kdjR
uP5m7lHa7t41qSsmtv+7wo+lzsEJHz5lafaBly13R4tcr6yHuNQyf8U85RcKxsIcUwwQKPfO8O1l
jfWRIazUXCwfoI1+DjcmtU9N4JUkvAbr6Typok5oTQCfHrojgzvPY0bzaHX2VhAuuEaCgV+a59cL
HxRRkyyhrr8emuMQUtx4QIn3dEOQ2qWjGR5heeJHM/8Ngt8vY/teftfRyjZucWKdTK6aCKfweLR+
ZrnwwzBjRuYB59w+arIV5CxMAqJSGls1dwtwLw5Pb2drr8caO7mXfGq71A6aImTuDPPL4csgO3pX
69MRL54oPNv45JO8GRdARF0DvkoTja8hjQmpxk4ZRx+h+Czdw2GJOm3duE6C6phdGKdA1B8ycuq3
ZJA7bP1oWoZoVT9bpcY9qipYrC5Alotvg0GM+N1g2cayCb/F2Nde2VoR0z87YIAETu6Wf1IsRvj4
gbCLkE/vHjJznwYu6ZBGZzzb6AJ0l8LplLuDfOdSL0YFoLt0iAlpPElrYa+wm7YoFPkV5RA7NxLG
+wDCnfmaB4bUBncHAjIktU883n5sMR3nb4VYUb5Nm6RGPxINE22Kn8cnhcmgqsNFkyhlXjP9ZLVq
cuw8toSPNWEpCGOqZ68cWQ/03WRDaXrqFbUizY+OigleFsm0ovmFC4wTpqH4Hl7vHr5m5E8a9lzQ
sqB0OsKp+QaJi2AyAF+UopcVxx64/pxM06WhEOC8hP3stL0utCW5JBRqf6mSHTD95CcW8S8dICZI
F2mSzJoCuChgTWkKhKEvOAAivM0IW3fr3mT/sgI26uZbgFBUNPATg8f++R59x4NRk4f603Xg219O
Fzpv9lopcwPQGdMWN7r9e/6WHyyb8ebvWNiZ2wuHH25WFFpjXS5eepaO55nq08rV55+sVABQFk+z
fOZNCCqDQpeHsfdW+s8KMiRBIW4dDHvbTFtHbLowR10m/NIazjCirY5OraFsByZAi1CgnjzzDlIC
Be6wW3lSQeT3ivGXYr678Km2ODVW+tI9P4MC42ziRMuDiC3sMuxHND6DWOZljHLOyjhj6vQTg0vO
uKbIjF+fkRSMAH4V7LmNWePVRzq/05BoC4CtpD2D8qFNbOC4n9d190nSYx2KFye2lrEERH1mYRQL
CH51/kz/8JLgYAlytSQcdbSsDgLPk6tP79q+5uj0zvQ2uu6wULWUmJfGo8hj9Yji/tJypnZ1ySmi
7wdoqafbzhy9ZvgQV5ddxc3zey71KH2kA5MUeaJX/ED4IWmGrl8YudxlTh3INEZW5VINC+nLWguW
HIJydhVdIg5XbbwTZySHWCVoJKrp3heUqHilKsNn4UG5DgtvXPHH3YwiNYlzpekwNFt+2A6riIMW
iBsgG+xNRM2sp3OnJP5uO0wcFtjZN98rfwOhYPUU0g2AxqZc1GeDmR/LxEGvVB59uMUIl9UzLOOu
qPqspGiIcE5abqZf4A4KmF/mYZnJJqo/f7zz0xUpW2MKOXlnqzwkjBErUYyVwCjzktbz/RhJpUAI
EdQxnGD/M+KBI4UQp7L2W6IGyeSYiEXt7jil+Co3M6xs/5WnQLQCSvTxZ4pZyy2EK4SZcOupFPZz
Mi3d4qH1bPf7NEqg3VzbXbBNE0QkOa+ZxYVOfAxpAKf+9/ExufYINN8Tg3luGExsRwEykYuHnFuo
5wthz/ZbQbywpoouPbZp4uT5yBj3WRNJmzSftBQOE6lL3ETqn7JmEfnmN/3KQFFTvkMqR7KZtCsI
NZaGaPNNM3Qyc+g3XmIP4f6V3LuOvvZ0E+pDgt5Iw5CjaMs3aYwkn1z+ELBWyPMxHX8rOVR5cCY3
MYB8YAIYlyDaw9U8+dudG2MDrZvWHPZukXqEDuXbTSQXP4lOp8xELvsIoSXEg3fUxmt5HMVVwNZ3
DJZfeSvLoQaK6PK4cVPZeziroH/57XP/aokhj/wm9ONBp5W9m8wDHZkq9FqJgyUlNbSnAJk1Ymps
3DCN1n/aY5rrSR2Z4fL2S8/KxbID5C2s+G0dhCMvOAk7gC38j8DRTOg4KgNGoe4z+HcEHxwDMHV0
4y1yw9XCWG6TDOaxGEMc3cM6h2FhytXyvyPXjizgX34l5apSb1Gm4awzHTDT4DYt/BAL1lS2t3am
nDMmCC9rkesxGM0I1w7xPl2MQJjiYRLVOgenQ14I4F2bAwNTV/KsLA1eQLULzRPFyFu6QOukL2vt
SjbQAGoq/e+uzIYwPodmQ2D7Z58Mnl/OuglJ/fdCGUWyknTsxoxp8fD1UsXi/B8cxTldyPnzhfCm
qy6NHOBDTcovCibDMsM2n7uvZWST184ZWmBg/7Mf1vRLAVzV/D6mlvhgYP4WwunuzPYhk0SQvTah
KZ8Df8Demdm5MpfTUFij/BnNIcVdcR114S5WxGeCH5dTIUbcVBti2hg+3KQBCRx2zdQnpK/oJ/7T
O4ryrHZZbitYQ6301ilce+0exoKfTTNui88S97+44F2pffqR3BELZ//UImcVzdaJAuQXhgI6PLif
WGeUkD/A11RoKJsn/kWKNefQvOUpNwTzS4h05pXJbPWcywHCqjT8t9gjZzzu0t7/86MMjzjrEKN1
/lV15mbHlZm+gRKSHAcnm2XExBcCF6Ys1TYC+kCRVwuYLhoGu3CeGc6Uc2UzwVgudu8A/ItvruwV
D2Lw4ELbQsXAo3/w7abZI88EXhgG/EV7TH9eVXzxItgP+7JaDMy7elQHPtfrzBgoNL6w3qkKOmQB
GjCmX7IjA4omFW7+qDJ7J8C2b4kujxnyU06BQqIIhB08NIzp/RpD32SMhuI8DoRHN8YBzkf8C7IU
CwF6feOCNnq3mhTNQNaoeg2ZN+mB2PpXpLQx3SGAo57d1bo8rQVi11MX/FdEj3GzilP2tIoZiBfw
ia6VnhxBiAz3gxha1/S/ItGxynE8Keq4nhfH2FQZK6SgJKNIQMqd7HwGZBhI7qdwroIIqJp+et6X
7q4TNYKaKBVTDwSlcaNmNM8sVPKOlWdDRkjg5aC2dHM6QzXKGsZ3eIcxOiPUI4u3GHU8W6amdqkL
17n7Ltlmxp2muAgAqUi70GEAK/p9sTr+A7LOZUGnetSL/aXlLA/FJ9Nq+b8qQo2jHO9CASjZP3df
pKueUairza0+J7t54fa34yM7tV+69V7RXGClis9xHID9FSpFWvZpMLMg1d6VUuIzPvM/VFh4eOC8
Lwz9mieA9ME51rLPAFgqPwbW7QMY5ACqhxRTwtxexkSrsbKBinMf0T97sCwEMdzhNUOmm4w+5BaN
vg3JErUH5Q+Yy88Oed2exXbGDFyxq8cmRlBeGpdxroYENFdbEasoVZZJU+Llm/0yvyCzFt5/ueDm
WFf7EEzwhRDfhWAm7qQrWJa2QpFdn70PtgSoyo9HDwZjMWc3xq7orj+3s1KRLRmbrghIqgZgwkWz
me1TQ8fQT9afdzBPsqxpObn/gE894g8o73zmZH4ZV2tuu0QV6pMCNYRvDOy8YCCbUlpeQRCc6BCp
xBoqVRSLM8jAP0ZKshFJVOBR/VZiUfYEnk5WKWHWBiRtrPIqTvfCiHe+++8iKpyTjY7fyB8bNFTM
gZBQ77/M1R8FhAwroFs2YnrbhBNto6tt+8nu4SQsEJk4i6RCV55BtC2735hdc9ndSos4ZtfKfaT2
lOk50ULsXxjs4gxFeWr6pHUC28QCKkRxzaPC8fgWgY530nHt/qSHaBIMPh2rNFQeQG9AS9plP1Uk
4MIey5yF4LuZujiTXkY2p09JF/Ael9v4J4Hjy1R03TPf6UNJcweJ+fb0ZxI+9nCHEHjv1J8vYGdd
O2gC9nb8reJ+c0AcFih/LSmeIFHe+7svs2pc9ymW5MVQXMv9az1VogtoR5XOHmeWQf/Tsfc+6kqq
utuJ6z70ATXarlUMbieBUMGQbKG0spIj19LoTqFrz+B7+xKH/tpZalXQVyuW6GNxofrVWsz7MwBE
aXKzs4jXYLQPvd4yXNWpPKv+t0Ls/5Si3mEAfsl+ZxhZPRUVqQC3IIs7LXHvk9sR4CyOBFuDZYZQ
HD1LaCiZ1hSOceywKmIdmPyYLnD8kpOoZVddaJAgzBEDbB7Pj7C7/8w3uzh02sVF5VY9Jn13pXkK
ChVEcXBumPR5DoLbELrnhbCjR66iuD375PVVpBw9r+c47c0/OImvLfP4TFLt7o/dkZbILNMCrf0r
Pa1/3ymbxyrKtIocc4sWfFi+8HKoeO/PP0HN5/Kc3TbdzsaqyClETgvq+LEEP1GrOiCHaTtl6O0S
XO47WdEHP7fbp1wtYLQon6JjFttHg15pjggp2nqqB3VJQvxTOsHPKL4pLs9ahw5OGLm4iVsA6pNp
IroPuBdNOWb1w56LfKkMDEvHTFV6eLLyONkEZ9w1yJdYieg1Mlv7bHzC4SOf7K5ux8V3P9KehqUh
Bb7SiSR3+BKkZ/y/AXFsNKbaYTVijhqPSgUHXYWUrBkXE8/k8NYMtpumx4nnKFgptdwit+6X2wgy
FvXZF21fyeb784f2uuvRvjgJyy2jGEEPcobUYUj+Jw517yA0wBpBldaalNYfRdQH5T3NfYKgSZhD
sn2yS4vMgnKel3LJWlSleuoMgAkPAJMS5PsZm6Dy+tSPnm6mhRkqZKkrztvQVHlYzTZhjsmQbyFh
PHVY3WYchYDNz6Lza1I4QbYfmQ3G8m2C4xv5enrgEeonUiKZwE8x4ev+Wl9HAFgfvQJczSAvtEvz
hTJ4teJJuf6oy2kxletdBBsmJ11vH0NdPEewkS57aVhmGql/YRiAcjGa7bxzkBaPwWNpLWEFZXkr
DNT+E4Wf82iTFVSGlodpBxcC8mql2JRhnDd4liNYIlnTD2KOcYmFHKli/vayWuzA0pFX9mREPkot
SuNtN1SLzYewZDwqkgUEKXYJP8a65Nk86vXDyp4i7dhl4R4QKq9QtC5hIcCQBUIyBdBaeFkS9FVO
IOgUIr+90xOwsZJwXvt1wV1blB6kLh+fmNi0c4BT6QaLYe+DTDzfRuI6AT8GCRUGCNSheNzSWPBo
rQhu8XEjoN0y9jmuBWdQXu6xDqM/igsqjAv6LZ3l5OJV8g/mE3iEVbZbIxxLsa2bVCiJ0rO0WVX8
UMZng/0DDaBgHPXj8NbRrdCoVTFHmJ9ONcbkra5zC2CsXn2/1hShLevjLexNuHBkL10VHSinyXJf
nTR4VlLmaFeEjBN+P6GH3R3log9P5nAC/XutOTP7sMmM9uBT/InLKeJVJWa0YcCBLl2Lf1c8GuYF
YtLS59aZowmp+yxTld/SYqI+XHwg+c9/OgzQHL33JVvNAWG5b/btG9Lx9e6lyLsO6aH47V/t9Srf
t4PpIHmXtvnGMeviHV1E+DodF/NO7756fI18uqEChCk4F6pH1/1vdspXhxoAu0ZYFu5e4BoNxUD1
Jbi5535dWEwF3g/Fezu5w72gy0RSRwqn8gMssqZQ0wz4S8GXJ4/NADH6Iz2YWcppSq8GDAL8QmY4
EV33mQB7xyda4+kaQMgYpCcXrmwCryxPSPsvquWVC5aVAUZYyyxN2r6ruMXPMsQ6/s65nJ1jrsif
V/OkSMxUwOW9tadw5x+PjfbFj70qrT6yLhA2knjOWLdDkng6Q6ndy/1XRlyJ536EdQ+LC1VL+LVL
1y08jWrEJmUfHKfrxDV24Vgy4mzD40HbXPVmTY7krS4d8gcNQ2A114xVj/bi8pCGFsPcMpBFj7dg
FBLmT6iRze14U0PW9PabYdLTIxK85NN50uuI5ua439cfrGLiSl9SkeuFutZxWPiKpYKpegJMB9+I
HlxuTIVp0bJIRPMUAZPKKi2vCxh7rzsAIL1q6kPEIIyC+ElwMAVoFuatpf6m4oZkS8busdYUZVAs
48a5i8SgG93JaW/qAan3JQTEi3lS1g+PwKcaPKLJmffXAmI7MU9EEl1LeWZ6pSjiL7TAxWbxp7yP
joj4P4at9nVtXBv+ZV+FoPSIrgz4J0hmyGPaw6o2AreVVXf9yX9gWQFAZ5tefj5lO0iZHRCVntZM
8IjAB5qQNoYfDnRTHwXjKCqSyqpqwCKEe35ihC4efXy+ffM0PquQ6g1pybva3xSL9SdvJbUkEkjN
yaAUXqmKu4fmUa4CcLG9TJXQ6Q7QlTdWkRcHHwpRtFos258gyR0e/hj+Q8Z+sHP+f/cmBxX6f/A5
dKIwiB19zTooxdvIbsGddDtxFDLhfF82pTlh48dQQnBVBbLHIjGUo7ATVSYrqfNGCikHnboO0k7/
UPowF9Qd0O0MASbOhDR7y2xSjpj6IRpILZAIoJhR/8aIw2E/xG/8wkyDbs+Yxs8J/wV6X+Lvs79+
DYce9yuqYvmdfHJpDqwra6GlsKG4QLdskM1t9hNPBh8bYBZ+YWmwLhABHSspzsmlau2ZGSSFMsfG
ncv26ZKfulniLQnGFUoL9PToJxKeLMv76ULSJT5wFdd3TXJhUH938XhF3HVAzhkdMVmKSc8dbqUs
y64XuK9IfRKsnDdvpuCkF/3LOJKDeFPL42q7a5tx6gAp6SYO/0C+fNJGaH7Xqz98/uoSeuQyvWik
KYVQawjwbWRJow1MvALjE+wjFTvQygc2xXidemCHV4OUEmTFi1FCVzBagIkQJqBM1I/WTCEO09H1
wOGX3sCQpAYDhzd3Ri0jkz2ZsrdADxm+R8PYVEYNtk9MBfLgxOCCRVp9gIvxJDshAnnf9FILQLX+
/qfOdG2EzGHLdWzYpZZ8P5X+ZpivF+ldWBcCbvF8WUu25mdEcGv0qGC+qx0SlvWYOxP86MgJTsDO
KJ+l+Xmjgk4cWpnsUBqPAwARG2H+TUMCnDyJG3d1L4H4uK0kS0X/UYkw3bqdU05iWWqV/RqYR35d
TC1zRmL/Mj1RJO1rpukbp29/ZiUSvtLjcPMOCmOjDJvwYv2NCyS17qd8+PW9iBEuwQS9cOSe9HGr
Fki9M3B8Z7Mm/EabDCfG9vAzqC9MLD1i2Qkdz4yG9/As25OrXjl0TcYzMLC0rveP/0cDq0twWjge
84sitVNA4u8M/wnU+cDgTiO2B+RbYY51Rk9aQmHwHqYhnaE6wcknF6riURX+wVD628vqYATOTGcL
r0mLkf3Rg4oeZPMG0IlnI/DRnwrZ8uxy9T0wJoO3LIPjeVXrRk45TSJplb5dvCJJzq2urzS4D4Tr
ywpP9A2FYhtz5cLunhW95IckwdhM25b46HSN2H0NxzaAbgqV54HxFkG1zPG0v68Xd1HYcFf77cOE
undU2Y2bA/pdNCb6Oiq/OhriyN3CDGYs8v8fXD3S2Hc4A+qQFd6Ac2HMagpKpAI/lfhEgQc7F+vq
r+HmjGUED+6swhMD7ZYIeyhAKeuw8uCoQZu2Xn6T6pgOQQsEIB/I/VEtvWKom49S0Z/DgdWNnC/H
0vy6jNMB9WHR+l/YG6Pslpbwi0y48qDCJyPFWNZcCWXm1cwcF0R5Dp/xY13aWE73bDPiPu1iZpqn
CM56CcjywlqLMKLZ2tb8DzWxKRWUgMhkScBCMlj7neguEzwRtwbrvH9qgxJWmG8FoiaZ5PvFMgRv
c9/36y5Pz8hRU2w5xfu+xz4iZm39u3CNVpRhppdB6Y2mlcPR9LY3BiilqWCqlC5RLb8iOYx7BFRp
BJ8LvC9sjdLYnW7M+enS2ah6TSNRpydyWyqKZFKzjQ+yBP31gJkPDHTQ+3OHscqdantPzpR4FVB5
xasiab8wB3izUrIbaW1CgrSfxPhTw4oGMyp5HXak1jX9Fs0qt3VjW+tTWia/IOEKL5ABZxAELqo+
h7gA1UALvhqIz4ynuNfLkErRyT1FfI+g1jRb7MvXnKVT8ZD6FhxZ3kOsOzbj10RNA95jur4ZIs2p
2lOKzMGjZlJ7SLUjyZBJYam4s8ujAsqYdRs/m8VOVTlLdOhaOeu7s9hkAO+PRcsNYIf979rKBj5M
h6fvocf7ndrCJmTSrhiZDEqpIO95YCYjZ2teZgNYm9nUsK+lL3i6MX7kzZrjFK/28dOlOku+Dy0g
Oj2WRMREQm3JCh7mCOmYCKMd+D0KdogiD+sOR7Pe9zD0E/spcMAoPzVBjZX0UdGs41S1zcUI9/jg
hchjCr/jfwFdAfVW5Sn/8j26/uuycbd3pHkmRO6FWtj3hNl4TGRUPlukQ5yIaadc+XOoKqCIDGaK
6roOgRxKGGCpSe16XPJrd/7Aja9evj/x+6lqH6nUH/Eu8nVV60C23b3RYG0S1UpFisNa56otIcA6
dWjC+ZDJOli9jqD0GMEBRdsBVavVTDO0WwJPkov9+ddwDH7i7rK7o+X60fJHqc0O3t0qxm4eIC/u
VlKerT05A3N+zaOxjdhZcvim40JjNywknhhy3LBAvSMXwNMjh2guq76nXofJeBzKYw66X1fJMFgW
Py10wdu06xyT0sZWXLleIyVx7upi/60J54a5V0akwDJZaNmJnW0+8Es+ZgWvUsTlw2mI7eFRwM+k
pKfGWfwcC9UNtH2L52AZfM+/dcobXZU4HIpwlPzau6nCk2wF0e7iA9Gz2IYO/4MTtUJVkvWlixvV
fRhbzE6Az9cHqEqra5h+7DrwmskKbyexiC5Ptgch/j5woyeqM3wzkyK+tmcxK+G+9GCmfx7zkh8w
01psTldWpge418gfYojG2gR/OPyKclAeVEyigQIYTHIH9jZcxYIfpjRB0Qz9LirzPQ2+I0W0LsmG
9uqpQTgcuNGqp6c9Bx1iaoNgJsWWi7PrcH2jWdPUuBFUfN4j23j8TFiKJtRchXHymjDpYWgFrv+G
MNn1WXxEo5nnoqbenPu4VlG+cok3Q9OAEKVkGlG+KYx4uU7XN2ElGtc47FdEkPpvzvTZEJFA+3oy
Z+cT09NWDtBu3CDWd37qycJNDoOp2Dv2ctqWBR8FnRjuLWwp6eXAnyAbo+hlPwD3ZZRQ2ohFwXg8
hn4d41/GBujBLKdBlLdh/haSlg8sOadvfxf648QiOinHIViDNS8vSxDmGHuIXd8a0c9YxEPmf91z
kJBm1ExljYgGr4wr0z6D1RjEvWOMUeummOGsNtewR+BkDUQBU+r8skNmWBJYIjSxOKFF/6nTpKqc
cu/c4LfAzuaoHJDtvK9YeCB0jF9z5jMUvler7l7wO98GOqAIx8LHDkSvI+ZdikIDEUDPP7IpyOzm
tiwLI5CXghWMG7zeS01qCV5WtF2ksx5D94dLP26ana+jiVyLj0oz6DHsjWyqp1TZhLkfOrGWyuOQ
mK52byrE2OrjJy1hT4zmnlviep9mGplyJ8JYdYkA6uICn0rbpRwBEgeX5TIwC+Pey7U8ayC55FQu
0EmiEzvugyFuIF0OvztSxWekutZ91+bpLBKuqkfISAiLYLCstIvziN/oLXbhhsEH7YS3JTEl94B5
FIhZSbDtAwFcOr4Kspnvpvl05K1OSDqu1S9EAE7jyxdmt3lxE7GfUFYJYOvS5YbqPJQ9BsFHFvF8
2YC4pCAl9nLNHIYJ0nOcV5dZntizkHUEBuSt0/4J6zh77GnGV03ODTNtH2q5Iqm00pSjs6mCARQ3
6HVUmIgbMcaRx0lbi/hA624sVflWVaRBxUi29OyWsU38lBkLMflRBa6DSeUag89mt/MMr8dg2HbS
/4pGg5FQBIZstbDc5TsKt38OIqza3cfybJFnMkOQxoCB0ZlraPuOl8xeqHCvZam2W27GuTkwFvWF
ym5m6/ZyY2nVknrmOzCBv0i2tgVp7HGKo/8aCSnt7PLrSYQzM3zbvUNJ6sf686PjAg6apFkjZHIl
SP5X7V6ABX9zYFUAWsuCpK7f1qOoYEwzeHkpjdG8LZpXcWLSkZdpD9TtRuU580Q/2Dau7heZl29G
M/I6fDQYdWD2M2u1K+qikFSRdS7BS4eO+q1NaJCNbBtcb7LpPemSQdgwepXwlzKAzTqm2lMWojfo
m0TsERD9Km7+Dd/NZE4wUVfi1LX+ogLMjOGU0eAu1Z9M5OoePWZiNJQjwh5a3InTzNFXECZFzE9U
CMIrj7F86nwwITZT8kdv1lrXvTr7MyluxNb+Zww3GAZInobkugsbAqMFHlU4oRKPO++VrjobTamf
PO3EYjtNN4Eqq7nz0Q/ziPwxJYmusaxBHlUZUzfOnClpHT9re5KgHN744qWIIdT9ctdM1mp50tE1
qPSZV8EHpeqhGHSArDT3BiBYh3oaX3NGCjyk0qsmFU+Zfb1QxDJYbJDfadhJ3O7JcX1k6k2VDI+k
YvnvbFcGQiCGkPjoYX/wSUoZnzJ1HrJpJIDkh2Zuql5T8WqvPmegWFBaTrCYX1AH3byIrUx7eThY
d10QcazB42JMLOX67xob9tRCEVD3d6ZYx0B29dUZZ0bSug9epIXMkL7RaopDGTClAsoDkTTRXubG
hQ8kPpT8HL3LiuQjzYRikm31/QjL6af/bZppYHgcCc5kZ3dqxN3YVz2rcBxRbAVr1a8Du5Cmvzpx
KBH6bCUB8//eZ19hWI2my76jmtnQ/cXJAsAYVpwBOB7AOqHUYyxX5StrUk41CIo6cIwzMYM8I39R
CdC3kWXVcuiuhVHhYfkrAt0pNyD8FF4FjzzdBAF17A86Q/FB6tkumJf71u2gNBOzb/fReM/7+/8H
5mvIgrrY2mNpXhVFWtHrqGEz8eTP69ZBEQIWtpQXdNRr7Z2EFrB/FMN+Z5szEIsGnZ6tq2MnLsyV
nPG6N5QrxGwwAC+p55Nxh9oEmdGjLA5DSaUYCLkjBe1/IoYhU/WJM8Z/HLFAU/qnbe9gwPOv7kJz
n7MQq1g3qewW0QjddlBsyDrWOqtJNjVfBg+qX3y+mY9njX2NpM6g6eIDEdi/kACC1UTvVZhCPaM1
a5BBhZ+q+pV93nxBdrGO6QTDVWkXmaskObNA1VFc5GoUTAePezSMpco+WV1U2NdlY1Z6a7pNs3cD
n+HicopybqK6aVqR32ID6InYDmPnbyOJbnqhCETa+yKjn+nvITnzrasKQutTQJwMC0FWRDjqLfrh
2JXzfEO1qv2gTAK7um5IyszmPXqot2RFrfXSaLi5t4YSylpE7rzczRJtpXaB6AsAdiVCD8x60Jxv
HvZQ2wdby/dKSson3aQ8YhTYBUSrmthDR1eJ5x4+VxWWNidhD7roWCk3ljan0cOXGq+xRWgf4NmR
sjGe9XhspICHJapXcTtGuDlOD6whO4gb/F8XsJF3tbnnQ7v3y6uijLSANlSwUbgT3L4U3+kPCrG9
23YPQkfAwYziwYRcaf/VbML+2SVMgFNSxfOr2BMMjvlASnIqJ+dcx/9Xp880795Q9uk+AZtLgfrI
Hvy2gSCjIt5/q8ejU77q2CJYkckpIQd/Ct15JmskM2BC6xqDeipcQ5Np5bHczpuMhZFpIO3Zzf5F
SI4yjnYG6P0QK/BszcGZwgnRUTqtSQHN7bJGV0HmR3mnxFtcSFzx6gb3xrdH2EJPsC1YGbBqwvqm
+/Zq15LTBRKJKGh5k/3JKxmUQzWtAkhLybyONvp3mTP4Dit/1HoHe1Lcn+TFXTRPcVURJMp2TyTz
VStxGaaNzfA1bWBB9zBLy+7eTyQ9w7JZn23lifIAB3dOWyOI13/bVzHDqqGsv3UhdXGZqFSopb5Q
wUGHVuDdyLPnkLqh6ctrMeb+bd+gH2jrU0y5YZFyH08me5EA9HMgHx4IojYzcZLU4iL26Bqu+mLu
+Ow+cNE9RNyOm4dKV4cgUvQWIzOliTfRh5jsZf6szqDn2uKPpK0Y5IUGpd0T/k5YSojSep93A791
SvkcT6n1S7QeDJHUoAotmpslzTuIMOJxYVbqyz6mtf31ILpXoJe3EKIEo4UJ6DYvswQmjIc9FWvk
SlPaOfvs59C6cxV5OerhbPnTpt05/CNFN2eJDEkVfk/Sa31NL0jA3qtD+PINnwvk5LWVmkY4SVld
41fEtqcufWYEMkUGaLLAKRxT/ripDBLskPxQ/InRRatA60IdDyVKUD+6hBFI3R6rS66sn1MDAojZ
2PHjSfwcocq7Qqa9zRhSI9bgKvWvxWbrcNspfRYRdqCAN0Zj011g7hQJtTAGaaYweRukE+Tqc/j0
RSuNnZAp8POPC0MUERkibzxP7IDae2rU+g3mE/arDmba9meH1WhUVah/rNf3kU6noYHk3eeF7Fza
qE3iS/NDQ9cRj2r4WnJj+G0yY51pONXAXSjHWbnsCxQz3MG+qa0QFcdSm/OHpP+s3axNhXZxpriR
XyfLTV0eJ+8qLDa6qQr9dpOXsdPR7lPQVyzdgfHj5mXhhG315Y6ljflKV93UiMp/TPPRGrpHTBuI
jvWJnDIQYBAolEBnvOfwYUmDq84ZS+3RQ/+m+HRVv4pdNvQX5mXLafXNMFicqcgpToaa6bdObHVC
Z7m2OeZhhg7N4bIsFf/L0cVj00mwI2bzS+kG5kXjj4u7dWN0qYvz6zbxkT7GdDOrL01ECnjhUwVE
Hi+//kSXsmO4l5ZLrmiFHxhlFXS+eIozn5O5yTvpg+BUkDMPe6KL7WJ9/NKa2Zf+R7p83T5TuCzg
cJjsvuAtVzoBPPTcFPpicGC8t5yzr2mrqzkb3LbSZb57EMxri4txVRCVPSvhTmCPyaDhCs1saL8g
AFNWyv4KWQyg0Biixk2bTHsAbr60mflSfgpSz+urLfSK7my6IvlZxEM4ddHH+y1V27OfKn8UTv9m
/jYcmZN1cTsjcCb+Tn1ZmKDfEeM9tK5caWVfy/2NjdOyMOAkCEk3rzDbDYAB8NPPHFxhuHpjumJc
Pmq7H3MihTUvFmPdWnBOGIX4FyKDvvcd38QZiTJGgNLrFhtW1UxMpAsY0G8cD3Ty3F2lOmsVCwuv
s+fxvHxhTLIm4gZN1oDfuaBQPHcQJPEecUlecDsgFnbfh6R7oJXoMqjjP+RS0DMzeWelTmSoeWwU
CLUk9NtvFyuluZNlH4tBCRCvtBdMjN4HL7Sh3dnzZyhulC6bk/+pu/5fUXAovgoj5Kt4FkvbF0wN
gP79ns7XkZhKVmAArgUY1af0v5kMcvnoOWnSPu2TLF7ZKgu0AKOST5q9d0QhfbHjHqainhD5ufyq
1V1WcG3QJgIFBEOZ6gda8N3anFYCf1oqF0N53G8y1ZoDX4vadEO2tegnoHPHM3CwrgaXH7ZSlL9e
A7uIimxqpW1AFfb5iQmMpnqTqUXbcHdT+2eSBruTjwdGQ9X1niI+QUYgaTmHI+m5rLXMXX+JhJGI
8ZrOQzU1QyIgDeS8m4Ts065o7dWgzd3hdFi+5Bv+N869Sx6v85bWYx445cqLe9xmOqotmuB4nDCA
QF5RQHkOrU2jYjfReYA6+thUEwSp6lJzddcxrqxqCAptXNAx5d+gRXugIuokv0Kforily1dJxz7l
wXJsI9X/Vr9n/1ztwXN3LbOJsdP+L9kjnoSuhbZsAKmPqkVrr/DNxUOQtXHvIjxTLkP/ECyCpup6
WJYEVCgQm/ko8Q1Xs+XPZMZTJhBCbLNSgoQsBVf7bG3dJJx55TCFdCLpWfg4m5jRrt1czj3NkBpj
FrinUxpf+GTtczWrLHbgE+9NCM2r8+vOCniDl4YWFUjMU+ibS5ybhpIJrnCTrgtk3VySIuD00NwM
m0q2hlwNtpKZYCOfS5N4WjVMxPwZ9aqot/nVOj45fCezJsMLy//1Yny1j1YHa+vBWVZ/ur+iCU8X
qYCfXuLKlnu5+ZvGvlHA7RDpHZx6l0W+5l/j4UhzmyIL6xlMxqZIp5RFXhyvxC/9S2SHBY3XYGFJ
zdVpxmY9vaOhBLuQXrVcSI+KqenYzmUu6TDLVfBraV+0NHdZAA7vX1V4hsqhofvfOh0XfbQk1a0i
3txh5M+gYwVhiH3XJX8NRxv6S5iWWg0UXCzMmXfv6Ov5omyJHgGgjMbXelL82LGHNnzgMIsoTrd9
TMl+jZp7pCmb3LO+ZbCXha2/WVuoaVdijQFPbl+vQDJWPvn1FDoJzqf4pYacSYd7xAdb6Yj4k15S
V+7MKXr6yHLjf0Mq9IUKSr3zsiC310WY8aC/FEJhLs+stwBcTDMB0qIyjiEiTioU8ssONacZXrSZ
5l+eWRGfUKaDqKBFUiV3y0gjxWts+RULomXbevfPat+Lm849kBId6OigGkl2Pqy2xME3CZ4Rk0KI
H+VDYaQ7u3M/BfGPjyprKScVKi6v22dj/NsMMNBviNVPMLsOIOmksl5p0T2uDHytjHWcaifQYlvo
Mw7VVQRpX/Uzsl/SMCslsQVJiXPQ4z+e6OQjeVtfg1zGpWYsudZ3UlQJZZFC6lu3MmLqxWJI2pXd
wKJSheitobsGbpfCElAKtTDNXsdrJzahwcyhkg64/LCd1gSXzT3T3uTVkr/ZGVjL/4T1GB3PyYWT
1GRkF3D+w4ul9BS7vKIIgEaEjkN+9O/vH53iXL0ZzmfwKO75n+m6nbA5MXpxC+1vXXsC1olAuOUi
xr2kfH/RIoNy1okKcdiTjzDOmH6yQXTp8xYSdjd3bTkflrN650QutN5khesQJnmWLdt6bObSMNLQ
D4bpvWiaBXXNznQqExEBemCNiGwmpTlsRhjlZlsZeuATfgeS0VMcX4MYzTkPP8DfW7wS4KwiaOVp
iyoJKxJjaf7sqWbElgWTNg8a6tF9pHe/I+E3vMExj2J+2G5HLIX+WGK9qwHQAjWyNDqI8h1g7R0b
RoK/riRBHY1+IHqmazE9Qd2X0xzp7t+kp+m9wjXi/6t6cK24U286W/lcNunOAtJnzNVTX/pe/q3I
BnvrFsRyonadG1d2Yd+1Lk1bDSxzJEwmOz3uBQkWgmjQP84DAqg6o2ZSEnI4YH3Emt7fIrD6BBnC
6sPp09UDFNscsoMRIt5GA6qOLGnd46J9bXa7LXvNIzwEyK1ZB/fHbKF7mVJVu4+0se35M+XzNJPM
LNjnegmMBR9ZRyzd1oFzHUgV9naF5IsQYcAJWSRQtAkfxnRKsqkeHrYMVlzyto4RMeFNBmE672QD
WjZEDt4zMknAhaaibAVwYoX5bGe17zLl1Mvp3ZpF+E20bKHRIMIyz0ZCc7o0QnquXuJlRMkqCTkO
oQSSP1TZhJj65KiU9hBAGQeoRWjxs2rAy13pekIvvov4vp7s7aVUV5dw2gwz2vcI4Ek9mchRvqWc
DFTtgt5nhEi77rPSbnOcKP42gftDhYRaqFW0wRWCcYWpcrOrMLcV6S03UiRXv0MQsQzgxIcI89D+
o12mBu0+FUWcMyAs8hxWeaA7FKUHlhPXF9h5kWJmCdx2G7MZO2L+X/oYohiu7x2D7mY1jktrtqu6
WTiPMJGmZLNnm1NZm/WRkRnerRuh/uNEJ6A7Kdi9Cb25VCZf1aH7whF/MkkBH4JeUo6omnDBpF1F
Z02m/dheHvr2cUmm4rf0VF0Rp1jtlNfAdOg9/SsxrT6uIpBX/cqTlV+y3k0H/rG92rf6ZfaGcJ8h
kNFp9f0Ph6l3A3ttkUj/A4hcHatSMDYExu5V1up3w3sLkXeWG574GBDjJQ21dRQKgva4kOEbGAFD
6xjtO+uRnZR9SphRdokUgi7A4a8J+mNcA4EO/LNTbNbku1p8YktXsfMzYmulrN7cGISSNyPlzt61
0GuYYfp61sIqMOkH6aif73x7EVXiJy706gDQEJvcuPmHQRkUuad/YBqk5/X2P8pwaUBNVljAjPyY
eANevS/ZD6Ou6na502M9bC8913qL5pZa4f6qVW0B0vkV/1tyeNH2dpfKIt47s5udfP6gH/sajgH+
T1rPIsqifIgtRusmx6T6HGu9e3eO+MjiDJTPI1KbVWWb1VafBwr5qWuOHdDhYMd2pu5JNe/YTlOf
LZlr20xAL+ncrcLrTAe2h83gwiEU0cys6ZUmu4p23lTSb7T+ESLRsrV+ylBXQh1NYIVRMFwZAT6m
6pQ4cA8wQw8he38vUF0zff4U6CdYKP89nLZIpx+ex55uCdcz+h8hAhKI5WY6Izz8qAsKyE1WG3Z3
OwduWcGGuhjbOv0ESJ4k8VSBQ6Jjkx8n3h1d5w0wOvSivxxNJT5zSxhmuJaGBYaKwBwgmtd63wUP
JB+wRd8HnTsCytGi/TiIf1KTV3rPu6hhWSaEdMNzfpjWRwOvjNihtyTqhzx9zJjIxrj7mxA8TIad
YDYC9g0B9flf0V6IBIeDnTqQlGo8lMewNWF3j8kNLwylsYMOcCswOewZ/Xjr9b8Jt2gcOBvNXAKf
Tiv4AuruNOTF6UhgNuRi5fRxPz7GlC/cEehcQ/2w+UGueVloFs5OlhVBpDQmle02NzkNf8SdmvzO
Sfkyg5o8ND4xg88ZwoF/k4RgAg239h0wNoPAWnOSk02x8U/ypXAP5UqDJtKtRnwTQsfOOQ4lYXSR
5MDU450T25e/5IDpSg1RO/HYqcixnmfcy99MzefbkFCsKu31d8OVq2Y9foT0+vTZbPcyWLIGqrzd
ewQzJdMdj1lSjW2wux30G6yuJ0Q7sLnjYbrYw+YoznmF6iPLjk6LGskM2vDEE+vfTRdARzz1lfZ1
9WG02iH9mnZsOBW3fcrz1pVlzvp3jqYf5uB5JMF5ko2Czp0aF1GZu+FdK7G0MOECojBc5dHHmFcu
s90G6TKA+oD8JuJ84mRAP9OGKH3zsoRfZDQxdJNuIelSr9ghCgl9hnVxeauJGlMUfu4SsdbVc/qp
u6SjNYJfUCHNwFxglwmzBlNKyEpWmk+zWu4+kYBtHSWBM6EUG+UX5nvgGIbDy2FvlMPoo5p5KP4k
H/+mEHqkMuyzyrxUc2VGLTL0QkbtsuhtF5Jewglwsn/3RefYzm6dyRSWxW4DoVa2Sox0zathdiaa
Gd5UNwLemycglSVM19sYyxtHlLGa1BayruQzfZdAYU1uQ04+L5uIFTdIilY/YoI5xXQ2SkIJeQ1F
mIpVwwtt54qMVn3nB2Lrr/iWMFUslQPzZDEZvoDzt0MCFTQthrwXKv8q/gZY0vCaim/lpdGykgaP
98cLOMFsfrBCBVFzDqvyD/BFGJD1Ef9uLLbDNicJiTMhpbel1nivNpzfoseKisrEp5NLJW8VfE9R
fF+WyYVEJZieOhrMua2Vt9njLNvN1O8BeDcFqYYXYvw7bUVhiauEFjl4LQlJ0OnsneBJDbb8aEOW
P5sYCjm1Q6xfxe+BjyVms690Wyvb4Rb1AgLEArtdSNX2aZd/BSQ9cxYdPacqAFAz2ZYB1jRjV63Z
HPVPig6oAQX6eTEIFh+m4JvugOaQCflD2X+71CmMqk/k7w6OMRLanFqeHNPXLfU4+ZN3W0eyjcUC
SHCt+nV3bx5V42G0qj5tvpOr0skT57bQx+1ZFek/+SsIDD1VHYSd6pEym7jdHwSV3+ErJSa19u0E
Wm8HkcpwMuclL31P0rPje4Ks19qtfFZq4UyVVM+9hDOF64d4EjVgRlucH+EMw4lvXFGO2ZHI7nVC
g5bNkn3FUD+5K+iYiZ2tyW7PoLRbFZDKR4NVl/7/6MiOgPdCyWUd1/zdR+5yTWd8sJ7sPRRRpw2V
2fOxlBA4c+qvtwTE5/eAbo65tgxhyJ6y4FOgvv18ulDswiwU+lMSUhX8oEcJKZenfKr81rUP3Gb5
gdE64vswLuf0ErnTAH+A/qxETa7kg4+TevNPFPDIccARJVFjP1bYfvJUvvxed33xgu4l2cqIxRCB
C/tKjjCYge3tIuycqIDCfKKfiOGAOFq8W9pCEQB2FhpkPB6jrMlugnsvDCXJ8xYShlHJkHFRQ2Oc
dVgroRd/GnuuXdKdAWvAyACxSgtokl/p6n52p7S3pz37fMQOcVBnAmPle/IxLQnqO7oDVJX31fJ3
zoRrLDfFU2Kovs0iGy28STW3JfY4OrdU7uFHSRNswLjMuNBcK3ZqrGcx/oFjQO7YE+ZaCzhu8fwE
3C8e3jTytJ/5Rko+qH/wrLTszPf8q9FDZxhFiuFhaCLxNuw8mENQ+UaIr1K+fkgk83iTsmgUq50A
3w4IvaXW9rKEQI83rJTY5bEKaQqS7o0nnpB76RgbjP7jUS+9NSXTkPvo7yiWywh5pgfr5C2eOisi
kptrq0gGYvjXtuOD8+5GDprbovaBS6dCLfE69vrDGYPWbOO6COl3qWM6sTKcIcfEUT9dxkg2Pb6J
nSEYF3+00XrHGLzb5CqTwZ1p0ZU8cvn6rTSJ5EGR2VRF9eAKDHgJtSFwdV81IaSVs/i6lG0shekb
l2LPVaG8xkJ0f3HlXovk218hBQY381VyEvtHY6Z4KvSm5ztuOrzGgbaGJqg5b2PWgCbU6Pd+XdiJ
zeFd02ynb45w2jXYb9gtS0gj0zt866THEbVOg9Fkovj2Tl3h2Jbn6A3FrJNMIfLhfocWY498n1iT
7h8m5cZKTKNwnD1XQ/+zwUnj5hyUJuqM7JvZYg1eohyQwXQ2DOHIjnV53GX6l93kJtGmYPUnQGhF
Dj53+9IzQFi1hgb9urgKdaxE60x/LY5DQVqOUpDY1cH7tSF/26yuALDYYdw2c8uuxLKA0C9HdiXj
am46D65Zv01SAnB1PoNRnxrlTYCH0NXbynZMm8+TpOggRoujuUB+BYAI+93jGcCamH2HKO1+TaYV
ys5C9Pr6TlwAqRnN1OeE52x4JyoihzS3qzosBRhfAZB5Jes1sdgWcbt1k5t2CcPA3rVeCF2LQJyR
706+bkR2OCRd9N2tM/Je/d8fD+2qBaAUastHiD9xPg/YOJcy4nc/Y0QZB1TdZRieme05YVAn1bDC
R+cGItHf6HrvqfAEgBT4CAJzBenI2T7svtLXbA7QzDLvNvxKIS0Ec2CAOj9fH4xA8aBp6Xc1HZS7
/sRW9EZD4mVbUskU/aOrXizVWNWg2XyluQtJfNcJgRdWEBa5L4mQOZh6HexxYaXM2Bm0UmjWaENV
LmyeljbYF52qcs90f4Lc46sVvj0lTAYXzJ6IOtyCWulMtFocshRoh5TucB/RoJO29ihtcfKt/O0I
aHdXWehOUrQQi1HLpRB5aHRqjdanIJFSkDtoRGmmoeWsKi8nABIfFMBLR//wnc4YpOjbDAuI8ODQ
kT6gPqTf7GRtDo2CO7xjr1WQiUEngIRLWm8QqujVpXDwvI/f9Q0C9qFyRpH77E8YdzHHXNCwYCmk
jwz/LMrLstYf1FNLaJTgZWIufCkSr5QKfGa66rO31b3/O54zbhWq99jv1dVqT8NR5x8T8RuCOyPu
RHXJ9oyz91dSL1WeYwBMpUDTSDMI3puk2gGrrjF+oXfcAKWvXnY+fKjhAFlLcp7tKThGKKj2YMKs
J4HPHYSUYHnnoDr6TqsO+VsBIwH0rEG/fbnBtJ7oIl7N/4j/xJOeP1Xq2qeieyEgmoRMVZ17qlF5
Mrw0CUcVBW+Rr/S2UbGIOnslRqYG7Rm/psY1OBZccigdE8FcSWsmKTpeuJpPr0wTNEA2XRV6TFVW
+op/spUrAU9IydSxleaqTpala1C2E/jtAnXRIMUZq5wEUEdKzXfjj0yc18WV7IKNgjqo4qkCuBu3
3nX5aLDqDAUqVbAwDan3lReRyUPtUtyB5cgARMEoR6mEL51MOEC1cYf85DG5yMCG9xNBeuaRzzfj
5e2YNhBxauQAqLGU2b+00KuinYZEXGuAcDsWVBzMqsNDAZYRULAvcxHKDxFALoAeJ+I4QLJH5XEt
YFO85chPL/Qc44pMs7OYeptWOoM0uCeSCzkP+A6VLc1OWmbp1DkBcq4nQSqjTSkSgrTbSm/7I2Na
50oqv0mptLF2mAIXOYxFeRef88pRYlP+EVqZqnYY5Ht6MuV1FNwGBzLlROuVZWDeEk3PNnp7vIsf
vGrnddAeVSf+e3sEje8lf9vooIxao9kL73UcIdojdxa1iqd8Liv561XiLwR2QTFSdsxtvTvTADJm
i1QCv/tby/c1OIpK6nbsrBPnuqxK5DxnHD5wCWEOldEoMRjM/Lp8J5Wir2VvP6aycIV9xJz5BkZG
iNPRXH4fuT2tjZYvX8xwX29xoV2WapxmuPeirAf0swAprw4dZybZPdrcoQfGrZFOWsfXNO2tW8wK
jokg9ChG2pDu85o1/onQlG30QtgBzLbMn5+dIyG+UznehsWcxIFG7E8HhxtE7F/Soy+3RCKu45NH
VOiNJ0+daAwFiugJ/dzPg81WnhZEi0/TTp3G4qR29/T6crsN+Y00Xi/eDHirI9rD4lk9MslZgOBn
hlbkoaV9n5n1qE1QvB2cI54m09lLvpbwpHlxfgJdCV04YyIC9ZJ9b3ADXiYwGPOnQuz/G+AMXZqi
/5AtUfxezOTPPblGzv/HyXI+xsexyhqEG6bNLDNe3/3XNBRR5AhUUKtfE0HZ9hGqC41vxs709Xbw
kjLU8KNT1mQ9uIFqba5NtsUqMDGMm4aecIp8KlAgeOO6xK8E8iRuYccyn5dNlQh0wTH2aRxbtn9M
LKQa1pVzfUq32H0+V8uxD4aFmrOQMJqYAMUvMu4m4pr3B299OAaLkeaqB0xEulow05B3fkZ1f1u/
Brv34PRKbli4IE5QGD9kwcA5RzgbrfmFtx8uW5WLeMKouf6/Tf8W8RzB+3r80Cd9A5IRihBcDuAv
te8nIRuUggdnXObkIMfbUYDlVEonhQcCTO5DREcdPttei49JkVmoBNv7Ls46bpGCXN8u9jwenn8z
sgQLVdRCQbGKFx1VazXeOP6vmesliw1C+tuN1n76FebfmnW+XNLYgT/9H/dOGoAviG+V0bsUHBoK
G/6nDTVD0d3gKfPfkRHB4bhCLcprp1RpM22AKwL0M2kFrN55fBVR3v0MYwZ2a24nhnxBaaj13sag
tv06hALMstvZl8yGmAKKiFBNwBmXbUpUXUeIg0SAm9lTrm/ZcUc69SR3gOSizHU7rms9b9qw0IQW
lw/LnQk7FHZ1jk/nPjAPMxtDCN8aUh2jGTUENKfYfwQErg8xhQIV1GZ9Pkl4yMwFJzDucfHauzX+
G3Ij/r1zeJa3XmQvaDqW0f+qxzT8mjnfGKaKSVSt4Xw6fEgL6K4B0E3iMF/r3WNUsKAVWDGEwQj2
KiLpRhuko01moSPL8+V7dyU6MIMoQvs4pogTLx8Lup/1qVHmJ/HCh2hs9AO55vwnucjMsGHAtDyM
PnhA+W9mVBFSR/IaG9LEVHGVEYpcFEqtjtAcBPU06xqwhl2Q9gX82csa/VK+GolCcUKmajXWDYGj
a+UpFzlelFSG/+KzwDCc4qRtfTjQHROd5ijLN0yCgtVsKZZ2yaVLF7/0viwD1A97eX9/japC12H2
1XSc9mR1m4DBU/8RJ1EuO2wOlnOB4evzl1xmlO4Q3kQxknoF1xcR3lGxbLBYBo6Ce3gmdLwkDPpp
+Hl/PN0b9M8MWZz04kiZujrkwQ4p5nGzEBOavJj0OQdhVZ+7OqG2DFcfvhSnBfBwz3mFP1+vPr1K
8MA0zIaByfqwEomKDPittD/mgYCRgJGU/rQPFbsAMvG640GP9fK34Kap/0mXioXMJDu75qpfX+ex
giK5DisR05mhX13rmQWW9J+R6+KEtMcc9IzhEHmnmZw12S8OZrxeOzSDMTfQ62H09DZLyPxatY0P
B0nS31Vme2trbRYCKYhqv9umgWyt1OoITxLB867RtN216O6QouqNyikze9eMs7TkLpYZgFM3bg6H
bnLDTO6biNK4c3TZDTXMtQ1gTjBg2CbQbMKXu0vB8floIw6ZSglJK3HUJfz0OYYrgb2W/9dD3fRj
vivU4ZMhhxAdtpJckyp+dttEHQXgVXET4dgP7xAl4JPMgt7u3MZQGCq1QazrFT6BI/WtoV+8tEO8
YWPyEjG0Qn9yRRyRpJr/igoWXvyM9iPwX2DA3cYeeSTZFSCZyd+UAykFD4qHevXGD+b/IVs8oL8c
+EEs/4Oe/WY8WODeMRMzl7jufm7ud3opiewt2TihgI9feUfNmzXmXdPXDYTuCXAO9pkCJqhLbd/Q
dAN1quicG71SFoR+4y/KNIiPuDhNbBkaA+3BHHzvgWBhFi1lHlaifRDiyOVBDs7wYLywtT84Jv9o
hnM2oZkGQohBuesuV2Ocq/2nt36NlHWkyIftbaZULTf5DBMnYmGNSWk4doJU9O9Ik5Yn8zQCyoyN
lD2jwUuscti89X0wGGuq09ayEMc5oEcnS8TniSHBSes/HUYucrWxhDnKwWiY2rzwLTPQVtsZXB0D
yilGpol07DqmrrFf63pif5+MxFK/rzKpu6UoFJSzsR/ygYJ9GN0hkJjXknaq9/WLS0nMzS9XniqV
i5+JO40sYPJY180GqI0zEJ2q6qV7i217TDlhyIaZm9Rxko9F7WTHJwXnmNoFO+s7tFjIQjssmRfE
l5ToBzTUybTpWm+ZUOKcx0NgSbI1rhQnb+H1lWz9Syts2+wg1O3Qqrn4BKfgCoImTefXyTk2hbrA
Bdd2uLdSFVAX5dGdSrfilMJwL8fxwO3B0LyjP2boqMxr3UIwWP3fa41xFSyCjKmbx8h9QU9pTbfs
2fv5XbvwXlKUTZ2/9R57ShOKTmOzSAk8JOHWhsuvZTZoTL6/X44/6M0XGnEN8OLr5ab6yQgzvzCj
141yYsy5ju9vcVrqovUipFHIAYtDuOLlGsqaJxSMsJ9UiU2r6yDa8I7b4HqDbDBluQ/1FDp9TN8W
kZQQEtTYG/eRGcXIq20e40WG6jgaAS86+S1CBgixxNeXmce/HzvRMSByjPqBu+ySB1ziSRSe4srC
8/4LPRUQaw6NC0el5NY0LnyOnUbhvlecqus638eIUXfNmrW6MVQvQ+SkhZ10e4CWXK+Sa0djySiZ
TEkVQgxhKaHKeTvJYdCyWAIZqf9XREkGVOh5yywjB6iL/Qmfq1CbxLrlQmzpO8MM/ZDLBnSQercR
wpIwpn3ww2demGuCvlMB7AF0/PHEwtIVnIQN3tLNxo0hEXaxiIaiSCXR15zPgKdN0kjNJizpMoQC
FrEAxw/l11I2WtInZtvxwWzj0iqkSP9htfqdCJiibEEI7Yw5TGD8D9WcEpLWHEe/jbZjx3rrccZ3
HWKTnRwZ2Wiu6OFpfwTJC8av3p2X6tUtG2Uacfwa50kN9SgevOTLK8GQ9Kk0dazEBRWewniRJk1n
GAp6GlYTLXU2sM8O6rrJHAvVlaYRIGxNDGnwNymAgichkfkZ4mm030gb2ZPr174K5JSTau8T2gKk
qeeAuBGqNRDITeKYSkaRhdCbqtwb7WFJch5N7FncszsERtz2NsyHxanh3zbiNnVoK3o7tRnONWiZ
n/pNcrCng+agnR2CtwBdeJXfuaTavIC1Bw0Y8BuWaiFk4c5WA87gz/Ji40o4E1H94t1HypS4MigK
LRWXNyCjqmyp++9xMazjK9F28TBYZ5NUkyBvxNMW9X4+Zt65uN8msHGgdOLgdUBjDwKDkZ3sr6SW
Hef7F/58Oxccb8QM/OT7ixwird0UGFVbMdF59KlxmaTFQidqXBtLC4TyedDyRi7nYBG2HHcjDP3M
qJ5YUdwlAQVpsp9wxKSfzkF+wY5vEOpaKdSzPOXyxDcj69gSrRq/GCBOWSiBnVzA7sCktXeJKIoB
NdRnM1tzPuwGDwMcWYcmrnP3rHdmbVvdU621Tv17kgAZM7T/MZqBwPO8j/0x1uHjsTzsyvzNHVDj
ew0YjbtHLE4xkzshuZT/9VjmHtO+wL6F9TBFVGjRT6z5EDAYIueMQhrrCZPyflWWKIKZtC6Rc3ZV
r2KqDUfsvPhaAgpJ+JXc9Jp0/xbShbbX/0LTPu8xhG8obhB9XJMKuk8N0ammDmbRvFcC+lryN6t1
U80wqa1ixv2dBDWfjzVAhDPxwAHD5ntlxMyw5OO9kFricQbJJ0iwpMUDpDSrwRJ86qC2T9fU+j+O
ee2dxgKMwCgVlsQ5z53KiJV/d3HuPIzBC7DIVoGhtb0LM5P0P1KY6OS15BtpMXh+cPBR0sQIgIFP
KEAXuqg2kiFN47gFVp6wtKrqIPrGwBYVINWZu254RWbeHjeEg22MWM3blNzRZuB9OyZ1EPzeHSYO
ODIrHpmE19c6q6pUQsLv1aPGv2GSA0MTmW9HhE2fxGAkT+YyG5iDTWPTWbNQ32mWOfkfYkmG1/bk
YkwSTHqYzKVCbA0tu4TUmH4kKet+OlZRYsnUcMpO5nozHqdLQ8KEVQPQeBS1xLhUqNBWRdzOdjvi
vGM4WTtacY64sZSNo+OnxpU2OL6uWy5uOQgbEG77HSlh5hcif8wJRSgM5KLo/pGnkejJzyF1wBD8
tb7/Gluxx2VscBOOnA2m0zgH1ChbpRGNgGPC7b73SbmYUWDB5GqwwerX3iRno8QExpwn2snuFYSE
W/xVb4K4EjRRdNza3L1Ubgr9tDraVjrm5TABz+4CkZX8PBvCEMrPkllE2ijii8D+Qo4GBG0UZa9c
b0tRgMo4Pkd1dGqBJqCXA7mOPedYU7r1965r1QWeONnavdLTNerIL05s5rS01gI89qtsjAuz8IXP
QsQtZhdWBpNFB7yN1gd3kHTDtffaFE9kbYEPQqH9+kXyi386vRudQx4VKlKCkBRCNbogwdY5zvh/
C+Jm436OiM5EzpZBSF8wexwNT0OXFAgHxbzHu2hz4OLIZMuV8bG9koIJ8otAPBLwQo+qxqXi2tni
EOOMKR2o42gIrJJUIlWzc/rjqYQqk/Fh5fY1D+ejZ9ydKgUIGNdXBY6Kscuzs1fYXJVINT2GcCbk
frQ99lIYzad/IKX0AiTh6TBfqQ3pbBqV8jMLvhKYPOxMo1ffPN1kZyeZmQpThzWlY5Kf470s5chs
x9RCJH5kIhc/8FsULr7doY4LTrtwXQEeMIUpxYG+rw8ops8gpLiNBBuSGhLRL9dFYfg1ID2GQx/E
+Ye1/RY7BjeQIp9Jz4k72ltV/COyhO/SOW63tk7bni3AztCTshBUbiDjtqfUOVwX0CxAhZoPKGKk
H8b3L2R1IdSG89dtPIZ+QjKmXOUeu09H658WxtAYe7iD5QVcBwhqi4gT5ZRQ0GtoIWm3Mmw4pWUR
JhCW/nMI6MvdDw659L7pJHT9xs670ta/mFE+q3uumkOjFKQvU7YYL3JFnNXjpQPW1V2FHvht3IbB
D6WsArvoZenW/WjhXIqVmOpNOxBWYL5+LlJbAyxBb2kRNFcXHouAh1p+6L74Fte+dFkB9cO4aoCo
aO3zvqho8l53ugYcHlZF6M4S1hQGMML/peChBIDEWuPhafuLj7voRIyO8DDqAyc8ows6xyoEuTwg
QOVISJB3mntl89kI9kLpFvAxkeQfPEcID+LaXozd6SaUycIzobsueDLKNS7lwa3Ahx+CaenVw6gt
SC48sQCtbU1191MYRfA2Y/ro37Oa/yOY22vHs9zY9oLT34JhatXLPztXG+GO/nH77oK32TnjRxml
xQotUnacZnl1Nx9Gxi0z2I/04GDHlu42y9+qEdQ/9JqxKtGdZO4UfuLbvhoOCqjYWL+g68uA4mYM
YM5WuDMf0kfCWbYH5vY8u8VuDjTLkyEjV03noay7BhNHMXEzKNTZAY3hJcPdJ/JJHnehcNkX63Dm
f6ta7uKng6tzQZFFJ5dmG6ERwcWw1q0/2Fah7YFmgnonSeNFWoFmlD5H4/lWlQdpwAxIh2zsbKWL
X4Nnbg/R8d+eJQfrFQa4j2Cbw0dEuPUtSj5eb5PqZ+GV892fJ4LaYLP9h3VHRzY96KmJjfGYRJE9
iaa7BGuDMzzzY1ZhddkmmVZpKmzMPcIcnf8js+gM6V6NHpU+5WjUBxeaZVEDWeKiawGN6eWVcGur
rIfS9prJWwVn6USFm3EhrBOynhZlARRiok9BWXLNkfLnm3Nd2K9EIU0uPsRKGmY4M1JOqU7KmJ+M
Q434esVwzEEjr9IS2Gs7yDLdvWXARjdJvz29jVAyOmjuuriIC3jH7qY6S7nTnB47P9pBCXixBdNd
f5keNXTwQ1khAj9AnpExsMXld3YqZ7vPCvJTmbWfMCW4LOo7Pq7L6duX9IDQVEg0TIPATdgNGm3c
cXkdPEUsBGe7B77/K2fMSMloln6BTFuVZU1i46T6I5P2rIgAYSP7MsoT7joapz4UlBYZeS9sVknM
B/b3l0lqRNvJiJ66TQeOmkPTju4lMhwJW01eTHghNIQ0TgTIadC68mzVfb6zBjsgg0OGVUcVLKjb
Bl0A2y23qHwr+zhxMEVdCXd4CUvPiHjb3TENtBWEEJjb7EFHQ6RSZJzRNWMq1gwpFQkbXbgR2Upb
h9Y+MhsfaH1CzHrJhIve4CzCoLkQJyOrqY+pPbZCn0kAJb8tlYlisLH8nHQuRHKHnTgElHlJKTv8
pMeAK9Ez3Zl5lx1bdwCgdfatay7vAxRftTX7ZEXMb9howhXQzbGXfz2Jmt8oQAa/7VcMftbr/CxV
Wui3X+n9seJfBVhoU/E/SN5VjcVS2Vdu4ZNI+1IegoeNN1UH4dGB4jGGzINql+hSoS+Cyutlkrkh
Nv4wijETg5MX/0wijWx0pKk/7bduFuoFY2Hr55nxjuot1Gr6wbQQsRm7mAMLqjZZVrE3THr0lUV1
4T/GVkA+MJPPP5arP7m3Gu1hBcBho7size8g/XAW4Oq8w8s6JG/EZlLqNoa6g9pJbpFIrzQLfQPX
i2+9Cw9F9xlzAg3TF47WkPbtRHXy8ZJyB2vfW/Y0BqNXc7Ba66sa99eG08ZVcVdV4K2PjdbHhhvD
W5cx4H+TQ+EgpF/jD6aKNBeMOd5No93ChY2tknLcPh+0gXh0DmzecRy51kRPNeSIKu58gvl419xz
y8pGKjxpCg1RFJbwHr+s3YwA+d90g13CTOiSF0AoGUstCgZGYrKTCygjCO7sFPOajAf5bC09i2p8
fFGsbYk1TaU43juHP2DL/b9xYNopyS6bkly7w1ibY9vFaoe84jaf0MojD8OJtWNTChq9fhOKKQgW
uURPIOeLSGVsDCe9FtIVDD4JHbex3iZz5UXkZywCJBeh5ywArvT9sh15655UVP7sg6NalGlsNeYr
BFA3DgsV0zRmKFEO5Jr27kAHQ9V6Ta36S0E5HqlUOqFTwu3EUxg5RUDZPh4Lga4a3ZmVqQZf7S9Q
C/Ccw4jiaLJ7BejyFVSWCNrUkCMQavyezB+0xQmVrvHGQ0611m2zEX3+Kn+nrikKTXUEolJe+61t
J8vPrYJEZzCmTFaKF8INg85vw19vftdTV+3j/mg0LOKe1758Jidj2SR6DghB8TRUijIXFZAFqjC4
+5vy5ov4q1qa3D6358P1wOGDq/r2VBR8gs1yqJuXPV3OwlHqr6kemxHtS0tcSI9mfHUOCGpvShZz
wiTBB3jiI/Un3OHLJCVWXa6xVMwuy2fuOBFhd2Z6ajjBw47Mhe9P2Yyw7d5s+vCQAYlkPOnlmRjs
dNzP2FJO+/G8xgNYtgzBbvhloAbAfa1rCu7MJPTQ1Kr0dfqOFF8+N2IUwiH4QZ/2moLcjSJ5n3Bf
eTrhHfKClP52139C0i+AFRw84kDida1iZE12tRHrPeHdliLsJZQP0w1aWDTuiN+R2mqECer+tIHP
4s0rcoHV6Y1Qyzu5LiGEbTx3TZhgj9QxI1ojAcI/pEPUB7A13i2wdILAMU8RNY7SCo824uutOIq2
1j6bhpgvOvu+q4Et3kmGy91a4FuaGuZ8GTyxwD689EnXylckEl6PAVqN+WdHcRpsNKBZiCP1ntIF
DpSkE1VX/CTi5pHJr3GmQUTTbfPQnQuL0A2DpDpR1MpmuUt9dLrnLS9kL2DsRBcfcZOxePn8EyY6
V2oeOh03W1muJKmWfAJ83mLwlqua2hEZo/oChfbjDoUGZxD3hFYIdQdTU5mAa3iuTx9nK9x4jjwy
vj1RqCnDbLbcqKfXlaYBrC7WLwOkyTQvq4cqcKi/+Zuc/xqO7dTVXzAtqeGGuLX7kg/knKAhWTfl
3RjY53Vo8z/9GCvdqIL9gCe7NqMTNZajv/2FMMbtJmO6QNmKGxDM9OI8UXdcIWWLg5fBUnduDzcX
hRO8jPpQZnXcBDd6l7fudtOje96QH5S3X656gqblJyMrLB77xZHpFn5RjycGXTc+eghQNxL8bP7z
5KESRVs6mLGvM/4xQqKMpm/639rgWf71rx2FNrc1OLNewhsmTTNl3xEll2huN8veiPxwIGsQ4/qD
MEomOVkuprquwUSJ7SqH4PumEONQ5ile0PtImq/GHYP2ELQMk/HslHunyXQ7RYQjk+QbBuDvG+mQ
ggybg6g1d8fZdXZntDDGs5qUEmug8v/rExxzYoUmkssXx9mEt7Mp9BtIbaxjZrM+zeL6feCKsEx0
v3/Z0TAAJ/V8GnrzT+DimIXhzG15sXzusBacAnd/wetuPBjbQwAPn/knjEj4gh3Aovy1kX9PNY/k
+dB9eN8lqjaQvfh50IWrQgCNkYKsZp1nIkvfEWj2kRuXIvdOwLddZd4DbV1NRJkdcx4z2I7s1Lit
py7ZOAOdOLuJxWWD38Ujyp6v2t49sNnhs0Q6BAUoRS9yY9YTynEjsL+k8PJNK0iN34RaMQoxx96C
fTTnEtFs8kzsDnX3kNJg8PCKroXUKQYqT+qZUfsmWYbP4YhTvC0TPRm4pXwoacsi3ZJyZVyESyH5
oVjJrtJyJlk7OawjRaDGJpkod2DwwC6jzOs96lmY4kl+wPa7TGyQy35CpXEAdKLN7xGnkz95ZYr4
REsHdqVZZ79NL02Ym04gPiADeGMcE+89GxdN0UBErc3xvvgHwkfUyCv3Cv3mRs1XijF/4Eo/ziA1
y/exv6IirpGcaMSUwAxEzB3Xx8a3EqhRVq2t2y9pQv3TF3/7rUcxCowFUfKfl2SZ7dGOXcB8ZYaZ
y3UGlAl6guah4+KgGUSy6bsKguWiVVNItSPxsGNTSLpTNFCzYXmWMVVz3l60MqsuPK+FMI7/MSqh
6tdYOmaoN6i62bR4SbyCt1v5jMkMc3bnKUa7UggF2b62qYeu7zSbxBrtAqkSJqdXMQ560d4DdSfQ
zC4w5fNHkEm8Zi/ZaFi5HnS5h7hwUV0Qswu/Z/l77ZCg1tTXDuS8nxAF5++X+u2+h2VQU9SqPXVp
Loq8U3py5KB04rZiltDySYiuy5VAyi7UrKcqOtH9HmKF6+Zp36bXs/QlKW84Tk1NG71KEWt2Rpy2
8oTtNdgPMEqAvmlh+dNa7dTiwn4Un2W9Odbm7qDx8cgEs5UUYUnNQIGM2qrJl1LQCaHUUO3WHZDa
LkFi201gclQuNVmMgtBGBA/d8URiCF92tUIKSTQjs52ZxIsrMm3Chq2/Tvi1VJTF4m560mmO3Vcl
a6KolNgqc4ygyeHNsUXwMBpqfoxLboeu1no3my2Nm1ytX9c5y/yLyAsXSdLWAGcXcUHXmHRpXLKk
9ggD2T33rbVZKyTZCW/yJK2ilu6n9PdD1JSTyh5fiFfOoUJiYaJnB7lu6NH1A6dZwGpoaNo6uOox
j3YqpR8JijWsYblLn2FmPooKh9L5KwypjHPZUej2Aq4VmWy8tD/pVHNWuEYo88X2kGIg76AUsx+3
iK+Zxi1Wg0PzunjKfjJ1CliE9TFKhGAABK1QXYT4uUHkmPPQHM4Donk6DUv2bI/cnSd6HSiyb67b
nwD7kx7IUUTpVEhJ+A6o0srZm5ZxDZQuGVcN3vl7J1PVs0z0Tn0PT98mOHRuAYpJ1gKYgdh65ptM
8B23F1afP4Xmx2SjW9VBa8G1VgjnDeFNLZo9ucmxPS1pSP0mE8ujg6VRPe39JJbHDsCoUe8Rqp6t
ZN+W7+5l+vi0aTVw+P1eEGbbgMHxMBVtsj+hDI/aeLXHKAAFRyYoNIiMhB/ROrCsI+iPR9oKH2bm
l466eqU3RV376nHwyU+jGsLxycclH6fpJ2KwzkZiLEbdTlYQRVepjwzIE7/WB95cxCtLlIMY1G3G
VkukVfeKK99/SWNNoklHwgHfOF9O91YIak4kbUrb7G5G0JZyuuK+QNsqcRDP3+wMq6NH2F1udpjX
DYvYoNhzzfPpyPJbVdIqushQ0o3Yh2yeFYAhNRYZm6ZZ/RlJRIQhLcIm7d9MnP5+RMKrClrNaKST
LE/GVCqXrwb/yFIxkmx10xVW6AvTiNotujjRin9zifWpK0XmnyBJ2Q0NfqAYsVMeU5pM2AcnAP8r
3fwH/swD/tmpQNcvch/DazKOwYzh3Gb5fWDEz00KGTT4yVUQ3GzsBxpa54YG54BDUxylypL6mehj
Frl055qxI2AjUNlxM9EVup74Gsr1P6Q60e5e1fhx0KrJvjVX69yOVSfGWXP4Ho11dj9Kf5uvjqcS
CHi2IFapB/JspeWBgAXwzM3WZvEUcCnz1OfFp7nETOwQfDyrl5whz9sIEpSb3l6XdqwsbJDO5wtj
e0lmnnTQDoViCDiSCHTEcrQX7TyqeFIsCTY1ksqe8hZe2EdSh5HzUDBpsNVfZlkAgaADxGL8lyAN
155HJCZlUSY23UgVA0h/1yvNdvUe2T4ozl7ahuMZ8yy9EHT8FO5Y5pm8xyUzV3SZVC0xORv/bOuK
apVInWXax/5JE/QHbzmDmCbMW6ZNnEZsdOJtck/zyImCWK904/GyOAv55155VPh4pi6Y5yGEoXa/
EA+LlIEfMDY66LrCB6gDLaGpsJ+WjNnPxs6gMbcSQCxbDHoDbXD17vm3UbtGeaeEOkzyH9HlFrcn
E26a8mw5TPzlx8RxO8Q6BCPK7LMESaS3vsPMGQRtnwK6MB8wy4qOffXY1gE0Hl+NS12DxBkShlJA
VvJO+plzzu/ED1OEyxU+/cplSBv5q+4GP8D2y+rTEWp+mWUbvTgag/IFyGQVYEAjb386pLo5GOKB
A0Fy0sMujdPBFtNe++JvMMfMq7ICDR6R5ctJ3S/CkKpA5VKokVMWPpwZAZ+9ptoCTdMHPEVG1bwC
eMxopPZ7LLgvK0qVtKGGmFODQQx6abWVkEeUceozaqbjxmAq9krJNvfP+YDv9D1XrBLCrQIg/SdQ
BHeqWNRDi4RB8n5PQ8GmEZabZvtbQ3sDAx6HZjDr6C9RuPVPNdGbO/Vg6+VXt5GICf2EGUM1wsWK
XXM9bsfpIBDQGI9M3+y0h2GlObN6C6om2HGwj2WyUoDCn7pa2ScRXvXoS4cC/SHmpdZ0RYvcu4jW
4dzMB8CyfbaJTVspEwKmHsMeNq+kZs7CWDl6ccuHLhaZUgx1NfJ+Hldnf31Z52G0UDQByCf4Qc/3
pcu2vKnTy6cJLo5KAirnit8H0/B+jX4qRY32kyrw22AJbtfM7AAPskvp1XZ2jxPDgsX+gZqndyBF
fdHiSzmRgLUtzZebmtB/x/cvsSw41Omt2ZCW7Glhls17cTtupU++WkSowch/Ygifso7jeL/n+y2c
y0vFMllpDFZ7FKFe8wdygP7MBp0rkg06DgOFP3koLoSU7kGqjWSqFeiZuO95qunFZT9rXCsPCPvL
HfNJJPhvnLrZzUYkUfNUQBBCpvUEixnD+f8j97af/d8OJCFnp59L6NghneT9ZwouSpZx0FT/Jf1g
bE2ESlbvTpkhACVbQGpIhautCEK8id0zuGC49Uve4jXZvqGdiNv6rN+n0rLdgPy1rxsht8Mas9my
qp4mBZtP7yI/63SO5MBHNBacsDgrFyf6oBCq95NpvLYEEBFEVh58BWyk7N9LEvaIDKU9yYO6Pt9F
eteMDF30CsWFaiNpxqsBkT1bwW1LYNintuZ6etDtrgUmDMuKIDI9RqoQoQ2y1XRIABJcCD1zoAs0
edyzCF4TBCfGTLCG4PBGKsHJiNVBuLzymEMag1c1JnPnKEjjdyFhnzr+Ekn9yEiRuXHLJ9Ih8IDw
lwj6c0gM9dQ/FPPcodpkT1+nitiUXepTNLUN+vEzU8frOpENKIZ7o2KqQ0a3s9uSY9QYTEPYfHhK
pSCxm7vysSR8JHaQohXcYA1Kk7wUu/Bo/IUlHaRewMXIr56CYph7xPLQ0WP7XdhtzQpAQMGzAFvO
i8xMFUd6LKe06h2Dw3sSVeP7YcplKsyfKEGr0wgMMM8gMivvs/AzY9XQBSql40YQjT55FaKfKpRK
vrpLWRZtXYueWkfudvE6nsPg+XvpOfPZVcWgz72REd4aeqq3oPpf54GhK0JeL09kxnBbJLOn0zuv
Thd8w1SfFfr3T+KLUy8D7X6ajcl933n9mXgQlbIBEvc5TLFd6e7arXUFDCtpXY50TzBDktKyq4JE
COR0e6UyPKLRxvHI29bcVmoQT+k42WhtNIzQIgFOqvQtEEJ26EwVmiiWiDtXbYuYprrUqDBZfpnE
SQZTccTl6soB/0UUoSwlJ3dj3VZ981CEOVfhovnbU9VBjTS4SJCfUvCk8f8Jhld8PTUkmZzVpIfn
mNU2Y3JUnCKpatCMqrfBi/dB4qoBoB30uU4dt2RDwbTBfqmB3JWfvNa1Y3aTEzzkObAUQQMQCLqK
//TMJKzh1IzbLdRaOL3aIiIM4tHke+6fbPEfYE9GcVkYuIVhvNeDC1roZhrCekYPEq7bLLOmkSeS
XMC+VvY5DdsGEnE2mtaPGeOYCKkBdPyD6zZKd4qhCwCva0mbdFT1dAYW7DGqgRqLaXHEc8klmIfx
Nb58/gAZ4gKe+JQHwJofVrBTXt5WHpNjWN+IjlUj269EeSc+nlxd0tnDXRJHOFQbSO3yaDL3Gez3
DLX9nDnmUM3RMkiBcBLUcI6qVDzkmQIsABhhwgAg8oj+24IRZAR0XBMXrCIrJk26g1U+jSOc+BJw
Eu2kzHn/2A6WG84lGpZdCH/n7AXItm5p7jgsKau8HyrQF92+IyaFUaFD9ZtOU5m1nWIQcjCblIia
XGIHsozw30C7Km+LpdiBQ2u0R/+KStL7KIiKeWRukpCiwmtpKMyLFOuYxIDcf9kqQsA6OaK4iLJZ
to7xnqhYnvZ5Dc5zxT/m2GKqAMwXIvQbawJOq7IJZe0qDFXQzOrszIX91XNwN79JKkBC/k5b6dcF
h8Ku7wZbO2GyrGvSBK1hvVj8mC4YhXsept+FSKs+duCD8MNd11eFqb8j5JJz59p1f85Jio2AUzhi
/jOiJj2yyrYzVrwrrokA7XcsLiWYpdOtqJG/jAXugcHQTKITAVuBsBN9/iQfi11QcxtLw4I0fPhf
PK1dIO05li954oD6FCZIIhbX8rTr53AQiIsYPRAH2xymh7XG4L69mTFruxHVdKsHodTqqdqZgN7v
uFsPxIQ+LnlSYotUlTvIufFazwLBLXivYbRPhbsuYndqdL4FUdq0sxp16Kk7PTSzZkE57pkAzX2K
5e2LvlpyKFrcStOtIOIkGYpxPlyHbDn28mrzsMiGd5SILlLWxnVNAoqq71cm+Ig4IoKCV9Eaj8q9
hQa26Ree4Hq1eL9MP49EJy6fKxsq9p0IEw1rE292TjQrFQl6WxvSBSalTgPGFI5U6Gm03dJzRkIZ
LWOwiKc/+0/SjjtmOEoAsDd9rwDf2cNU8Q3j9cD1QrLVgfywFNxrKdFUGAvbjfRiCrRK+NFBx5zl
TrzldFxSzNFt0ZT/V08wl4wUXW4QI392/45HFFZGB0s/Y60M9SkY5JngB7BssTVusYtRWmKj0IHb
tv0fz2jNF+Hv6EbdcTy8tiQD6yqZokKq/IaNIrGaXvZ8eXj1VKh9PE0kkyMx6B1V2MnX4YbmLJHr
hLxFRp3Yaj3qHWXFgyJQj2S9+tU27oqr7/PTpoeGFZBq/6ytbTwHyjTzR8E+teOS27rhTZokW5l+
F/8Lr5DGpqWvDKnnw5KhIDtHEj5IPt85ycrSs71KDdkfXNM8BX0KeCdVLKwQ48+NXv/00kd2/4tb
RlqyGY5KMlzn9towlu1MaxuDrlLmTHKVn/Xyl4ZZXchZEvaHGeLWUEpX8kmuMqQjm7s0CHlFYk/8
j313aBGN1sBA8W0i/VaojuYgDLYEx0UKKR69ImeqO9SSJbpmgTj6fhigXzX1KHX2PgCd0SHHW5xJ
ejBOL974/kb93IdReoDYtj/399MeRZkTIRIwZpj+bRKRGppFAHEUTK6y/XHbKxTw3kUFaBIJGLBM
5/mpeJ66qEK0N63zwlla8Tva/lpA6E4+pTNdYSxAyowtxyLAbmCruJISsRa9/uBq1HVdFkgs/eU2
uODIsHvoxhBhVwO6q7WVLdoRsQcGI0XiARvo1jNhjlQimxxpYFNJT7cAtgn/wnDZN04MEYrcj5zO
bfVI5MRRte11TcWnHpAd2joWKGd+SxIfvRSBhkATDoNluoRBLkYSx2iAEYP/VGp+pfNwoOj6H/N/
npXiKbCq1NqTYrT9WFboBbtXDugIkXYkvEkAF2UacqfbW5JUTotB2qsbNMpJkI/BPMBv+x2UGN+u
d00xoMK8lS+Q5WWtKReKYGUytswD7hsPHP9uhoEJ9WBn8Zd6cwEplfkLuXoCiigbHfqYUFA0ZQ2Y
EIBS5xcAumvlNUiHgJMenNZKijYPmzCe116jf9NO3CTEOPZLUE9fYTq5HAlJrrfg+QYwxaUxc2pJ
YkVw6BKM496TDqTwGr4FkZ4speN/4287kUPPRZH/iXARwgFygzdnpUTw4EMMlEdbEQIazMjyCaEl
mF9FdZCf2akLTpQqB37Pdnz51pyJzfYvJ159rHpOfw/pkXD587lFkjbJt58028QvTN5n/QEF7EaK
kq2G5QtiwTY3HjeCVtnJlF6ew7s9fNSg873Z/Sx1y7gptyVzgdEsixvyfWCVOxLoELxwjmAVmMAP
WtE3CUEvTGMBpsuR4IBdCuaEi1Ar4lAsK3xIBejMreekSqyTk3nzV/zw7cjuvnhoGJP6rSMKXdd/
OntGhYY6Zl5t5k/OaAAmJRJs2r7j5xWyPO+NonN5M4qdGMgqNsLBILDbmt0zLa2P2AKPN7p3fzkw
ELZUzAYrLbKdlufO5oF7d24vRl4egVSeq2X5AFCm3sfao7y1MOVTKF4/m2j65nTssZqMApc3plG/
vTxReXCNlYnvRMXi2X4LZ2tykgd5nyz79YHiNMM8qVev3PViEk3n9roiHwFJYgffPGh2CB4OhVGz
l4wMEZNeuKmHS2cmllMwWz73NYyP/mYodj/7OU24UgbwnoFCgVPVUh9fWAqpl66e2j4Zk0Oi3UXb
KsHem6eV/loEDaAkTNuHtvrrVTx6sEd5/1d5K+l58Qz6s7tzkPfha3JUNmUyt21XNYnlaz3+2XRe
T96pyciXd4oZe1LkJsMgoqJ2Tw4DNX2lVQ1K7QD5iibwyxfRav9Ys8+PbCYXqCzUw68LgkZ2w1gQ
uyqnkowv9UKakcYIYRdbosjhXrDVmGArWF386CVZ2hslG1c3t284s8pYa0k1rnpiwqoIkQGGIXkM
GR5PmGIRrBX7dIAQZCCw4WnqW2tN/eZ2hqv6tJNbG27lgAKR0jhAAYmH0sLfE2ptHQjv7uLoVOJg
58QMFdJZ5dna9GeUSP5He4VS2VAEphOhrcGx5PcXAdUiwEQ7ws3AGaOhIJZpjvQTTQUqqFNc6fHu
p/rdm+mDQRQBlZJrf7Dy7LDR9j2AAVhSzcsw31CPP53uinuZxNx81P78DO+qlnpXt2UxhiODeXDO
7dlLUGUiUa8pDiG8vsQ7kNvXFrcPIpUMv8B+HW0nHImDAa85NgE97elhO85E6Cx4H7ZbscXcHs5T
5/FhEEuLr5d1ocNW74tLk/3ufqG3wWaxOACgoqzNyW6ErYGV3RHkH/lWO1CedvufMN9OUCpSu8yq
sZf2eu7b+N09t6pidnzfo0cIiiPmVr7x9RkC29k/ckTmRBX4yJcvcbPbmTE0dZd1NXJpqkJ061FL
gpFDGVN2JT+GN6pMiVTyoQG3okZAu8OqrO1Jg8oLMFckWIKfYJueaJ7IiHNhx7BOHBK+f723kC8Y
3wN/JGbhF1Q6FWWDI3JXtrB8V6xR6LmMm1OXV3xCIJwsNlKCHG6biF6kj6v8236t214L259Hxw7s
aA5BhKxCfPqCdGZAUiGcmjaqJKd9lpm58PsDKYxrxaYV/IvTbt3mUxbcPLd9EY0FGD98mSEt2CdD
oEoW/mphrfs2ebKQYeXcOitRHIuw1QnZmw71VEAiW8Dt4KzggJGloJxyBq1cswuB1p/TynfUroPu
xbzIc3bNjFBEApnJrwdkpMyWNNvlbPRLOKERE6JOpML3pkqajvyz8t6keC/x1TsxsbETf8Excz57
dVkx1dOlMo9A7ZRjKWr2vxaO/tGansP7+tZM+N0KCm7lNVi75H0x1zU6bXwsccoptbDm8hr3Qrpc
Mbj7POa/8130DJ6AzZWB9LimOv2QIczaY3D7/8+o2L515JkkpyDH0bqJ+Jmnf9fmh2vebhSwGmXt
r+kQVTh5arYvIBvD3EYiT6Fsp4ShU9l75yPo3qvDnbcbpV3uuclEeX78ioILcKiQoo8GVYpjDxJE
Cc7/lIFcDzJI/44UF4iHuZ9aP1MOVHaF1xPKY2RbX+wgb41kCprLkChPQPQePv9SWlsl+JQ4/5tV
qLZ0MK5nCnciQCPfMlxhkyAjL1UE1hV/wSDGJtDuX3ZA83fdV/J3haqC3lqIhLnefmrmk4iubNNU
iVxDt+ArvODyLNskgMdZEvqHlbB+LOQy5tt8o68SUG33X4ngvl0MRklcHp/5ZOHylRI4yVCQ47rl
LY0S+CBHK2MREVXxNTI5W9sIJBwcLO+njOUY3iQn3wBEjM3BWzqkYpZvj9/P+B7NjQR9OERnnUqT
qFaF1KzvVLN0wKmhiie5h2DAPznhF0cFA+pYsFV5N5YqHUgOuD5XZTvi6XUMOjUtVkfaEZm1cPz2
u9QZlyBdo/Tg7MMsJL3o8Lx/JdAXycq+CZjbePLamPWvPDD9lbnpayR/ASepNk1/TgDnwsNDUpe0
xIvxfvHvQoHHUMDssFmHGb3eBXkNuBu+NLzr85mdyiVRZaBmB++dkAJJZbrZeWstSgSCTQ+3hf8j
PnhUboV6e/BYQysS/UZxBQgtLaFkHkLJHfXD4PF1cnH2IZYWDGTB+q4Hosa8nbEhjEGsW6Rhk/lm
Vm5ZtVcezmwA7LgrR35rBuA+3dHcKUEd85rWu2MxHgmRB9yBYQsWhmvjfWbDjBv5rbaLPFb3YOQv
UQc6DRFOlSK+ixm7hbiQl710szkv6oUKn4mMhQcinfCssiqQ5ZofK2FMhzNtIryw5CiMoqgcUp6m
FIyHi4PV11wXQtuJ5rPCt8Z+h87mzfc2/D56bhj4I+ACWia051DzlnXAlc91klNkcu/p+5oAZyLl
2mgt5sYviR2jlC9rNHV1Vh4Zx/hXSN61mEzazkH9rZqrE8bpghIqF4RGgO/zPhycgHhWRSZnKOKE
lpX5IIcMnykA4wr0mHFcTss1trE0RESqmkqa43vkIa5gKVna5rSoH/S9M2ZyCiHMaHy2ZbVPujuV
Ab8J+8VzHf6WAvIv/tdD05TraI+aEG4C30pzi+eWCgEs+385Op8xo4t5Jp0CtGgux4usOgERB9HZ
GsVI8Vrh2tBQoIK+LCOHzABT+zZNYg/3FCmrOVqLGifW3IOqz6fg+Qe+BPdA1rEvnERLQROXJ16G
nTzTvnU3djJf8hZHecOhtRTIIfcGOYQqZtasUfC5DEbzgz3Vs2wpaQh+tpqxU3ijkFJtDLy3npM6
IqBA4mLPvg7pPm/q1G65hubbySbtFYqXzep2EHFYnmiwXtBEXHJpR+LPCTlI6sk4lkhNahCx8MF1
OcgxrHgfGQUAbwaVk0dHkyoNFARybtrCVcqBZT1ET1PRsjRz7u8+MEIzdX0uJLf/rfqBTJni7coC
9naxY7Ke9SFeilPZYEMKjEAtiHh52EbXAJmgf8ylnpK4jeaifmrHwHuGUzCMxcq8NkudFGPRoxMS
Q1nAbvABNa8I82QP2hGxU2wJKkI7ulB8DZnwsJ6NWYjE3w/88kdSdAM8VhgE2SEdZ+ZOB1RMnJ+A
+Mo5OLbYlENSivOq6JRFS57t/65K0A8ntqRkFpumzhBw9NkTzTOHQItX3ijJalX3EVkQFT7BIhNw
iXTm3hrxcjgY4rclvxr6JjIt74fkFidDGYUuT5E5bBtXehUB5vicNg/y0kIwOpHqzZcZcv1NuGnS
YXx3q59YhpcyDDJxNVM/gsaMICXGmoJGUioBYTWGuVdR9tUUDdoQ82fmdpUYV1uhpf4W+rveJzl2
+uPL/+zQebJysh2m0zd+SXEeklM7B0edh4GHNl+7QMF0dGM5rcxJL45M4ncT0PmLaH+SVhqV/KeJ
9iJljfKApBFwmPmLda7uFofhnkDDkyZz1xAeyav2nMQlegsskZPP/5sUuSfSMFRG0WDtRMCc6wYo
yHwjHpmYpbtsj6UOCR79N6+bjEdXQ3ND0Hb1y8uu+pH94a9BDA0Kt/PWox0jKpP9XymdoB80hz2D
tUG4Y2xosYYqC5AHLjWKRYHLqa7Ygs9OUivVvCNzlXxkHSYpFG75vPMSlKxfXX/KsLB4CzBu3gqL
Z9I/ERiAWBsdYpLUBYNpqhYqnSLV+cYNCg5VpkofSL3g1MskuYj6XqpqQrQbsyaeC1JeQuK+P6jw
NX50M86cuzQmcCVItWcpN5muVkhQUicY+AGLzZM9dPT2F4pg02iDnuEdipmow7v/G0/it+esymEa
ZenUZIWnXAomBCiAFieSKEgPU5Jl82dbfEre1kQF8C/eyRuO2CYMMgM2vCPw7h5KW1VVVlgwzMiV
/K0dm24dxJ34xWze9y8oxEnFPgbK00fxUglSscruYs2jgkWlyeSYBK/KTAGzP8w2uqLgaDB9jJHH
saywyyT/MahOgml9wlwA4hw30iODw/ULQh+KaQ09zaKcnQbYWNyZBYCfN5O/9xBTyQt/oR+Cy+Z6
Fj1zWEkePrCp4ZgJVMGRXYL8YQC6DOhPqYhsEavUcZ3SIusq2oupWdMGrGQb/BRqtJzFAXzgWoUS
drS+3ZAHdwE5xNi5i+ehmIc+Zfxr2m/1lbZmTARin9R26iFxGFePGIAliWJT069sYbagRlGRbr3E
4/Vww7+JAC1s/htU/ZS32hXINiEi6BEk1ZkpdY+Fh7KdTF3ATGkHe1Qxo/JyU7jXvlxsZEoI+IX8
uxYmCQopJtUNHgFx/g4i54geOt1j8XuFsFygTmJZqeh4X5QQWZPF/1IWb2HGrUNQRRdy6DXca4uY
Ru85Q8Mvadk/X7GWfVVjKgOWJBKHX1mHranWIngkAl5v+y5RPlbGzEP8qZ0kaTLdcBChF5EyqThi
y+QAY9vwtaxOniRPmORtH208zx3lMdgst5cY6PWI/apMMPUZzMx0TDMLXlvzeLdJwqCh4NAjBv0O
+g9D/twYN9MVuUtZW1L+RNUjHpbUz+eavcVXygzg+EqDhpEsQlyYzILE1jvhgrHmhCoKtDcSzpJs
zQI26a6FrslAPjKmXhVrKUpWnpNOYXo6Mh2PKblVUzpKeW/vn0OPrVm3O1U+C+ykUUWlr2Am8saZ
wtujj0/NIT9tyV/ksHz/iis8zBrnI5YJ5+cQrfbhXFydHTUN/RSjnhnB7+u7mpMMJFPTNxddHDXn
zd2gPo/jdD//adezrB5R3AiFafRzVJ2+GnocN+tIhnwLz5HRxBNp5UVYUd9wQ/27AlRCDHHzcpzr
GycC5R7dHAAOUB8LOoyR9hHwUqeyDPyW++HHJC/9vL4rfZf7xIMfOcH8EbA9zXd6ZU3a7yVReIdp
SbO/Na6iD4vXxFCENN791nHzuauno9IETLiFIcnTXJqyHhyyJD8P48xWwfdFvsFmud3goAI+XqOA
UZzsC60WoEljh5xD3wX37xmVJa5gI5B5PY3HJy638gCL0F5Jd4kX7BxWShhpSENZCBaC0PlhoR9W
NazOkiHQsAyo/b4O181FDs5yu3DjQHJB9fCKNGlVdFwVAia9SnRbjc+ZjwudYjgaEKyqpHErXj6/
sX2ri2kwhos1foG3grHXEPTnhC0MTMflRu33SFi6OzHSPh1k9XEXunqI/U4AMm9ha+WlkwfN4Dw+
hrBEJKG9nmSN9LfCTR12Qrxe+/n0A2f88pw6QExtIxSvjnym/v68yBxR3V2ZR3Quf5eLu61TRl3t
/IvYy99Ny9bnOweEDGRgV23zCqW5YO1nH8Uq5dHljs/4j1ToO5DVTPZMegMRDkWXEmHiIRueHTMa
JahwNOcE3ZbRWMxCZMISOKgpFmV6NgcFtalbQ1InAuW0FrS6CUVX4RBnca/C5p34GWh45S9CEJ+N
R/XJzaGwkzbCVLHDMxBWzTQAxEZbSa5995/pG6PRoU+ua+amh3oDAIGgCUjkeC3hHC/Pa6toI271
epY7fld4R/VtVKiNEGcTgefbvV6u4uYm35NrX2ga+cM73luyeo1TMpGZ4c2A3FHU79C6+RSEy++7
auhQEgb5NUGc+CpXD1jDhAWSXOIx4YQNtcq5P/1TmYjC8RZWn+gl13qT9NOAR/HWL6pU60QvH/Tf
Tq5seSbkCD5uK+gmM31vSvdIuZn/iwDOeLiHxxsnUvPU+SLhnihdQpWY7Vxt2I2NLAU+J8bYwufP
kveGciCNtM9cvFdpmQgj3Rx3cDmQN8+PsaDXgIjk1P5tntMOjdUOwBQUcxQSeXCgQoqqA1WMPIrh
x1AandnNAqPyO6gXFp4lHKcaGN94NKwvYl+WI8JUP09pZW/6qqCMOKNVC8w8tvaZAtKVwFIE8KOq
I7ouImswMcobxHdKfRd+2mO/Vb1BTKEnfIZqcD+NVaDncsdA4k+CzIpsnAdwtV+YA1Xb0vZl6QPV
ti2dhe29TiimPMlUNiOlUpWj7jrXlg1JPtmGT3Ef2N7umITcPnEKmbiSUy+fprlZ5iKk3WHWHli3
WSPjP9WUisr6R+tQf0wp5pj+8lgFLXjeolc00rPpWhlMCfygyq/JrPKqr6q3xG9UGa5j1DQhRs6y
wTJxl0oA+baedVUS05v6lrMeNJdI+Y99WaBdqbybMl8si/EpX87F4RmhTAwQxEQyl8XdLLmxuSvz
NCNLfRRKPWAIhLHXkhmE3nPDiyVp0/5Ldo2CvNa9AzTWQRF+N0x0aqjFf/lXGltb2e/FH4nDt+DQ
Ki81tKpQeWSs+fcFaFksEFFRCOaud1/5KfuVdJBLcIb2VQdSa/TBKsoS2hULeXx6MEbUeph/ULKg
8kMHxkVC5Rur1QUUZJzuFatBCbiK4lzQVImg2kiMMjwVtCHxOHHDGwt4xU+E/daGi3naDxm5x1va
bfd9+idmlJJoWTe1nisLdGj11QDh49gSJej4G+suwRoskSy7eGuH2UQpJ5ffl7tN1s+6LszhiNrh
X01B3moa78LoMlJD2bYJ6pwXCL9MQf1xZA2dDlWEnzDnZhvITEkDATJpke/vp2FJeTXkZmWfatlY
qfTPm0z6lOx1bRMllbpAHLa2zxDrBpQF3+jWzoxzYLp4jD7ltGA0n6bPjANEyoHk5vknucfzThGg
EMipWeWoiufqC5dkuHxrmJcGLmWLB27t0Jb81Yb50l5ZILULMaifttgyhGBlieA9EkpJLzZLSf4N
8ZiWREhQZe6rOrVDKSEh1a2LM6YuJIDsyFza7QEGP02DwMu/eITkXlqwEQzSV67E0ti3UoOAiz5O
Prc1POP1jBO6khgAnaPoxvwDXLdPDb8EWabVgPvrHFCEcHcEzCTKGlDBbL7KGWmxu5Vxq8lwSjTt
iwynmKCfgyTo0AUWYjtk+bFBH5cWwAzUOVtC8GFmuf40Kmgp2XlAtyGX+Ugrw8PCBpzJD46AgJS7
elOj+TzheUfLoEN7hGK0Rql0lMBuhH+8y21eNNj8bp2poMuAHKD6QZgY9ZmHZz+Stb0pECc+FzIc
F30Ev8qOT6BSGQwHwt/pxiwdsrseRNxWofmXN3Y/GuMZjVjerTsMsY7HiZF7GH19iaS2OrrOG4om
dg1owJvbmNDJ/QUoSGuJV4DyGuyrpaxWUj4HmyCNylP5SenwDxOmH4InA1hoiQ0zsIQ+vyfxEoqa
G5QgNvP2RK2Vg5GUHCM6fl4/451Vz856Vl/4AJ1W2GDjehKsGIxXQ741wfPklJr6MEHNwcER43L6
D4lXLXb62DN3M7JRb2MXkVCV6wtDEfs6Tvi+l/5VpeVA3LK668VbbdP7pS75ANIRfO858rNFmehN
xF2+pK0fw4goPsvTgS2uBF2oac5iU4lEQOWybuBLqa1BvLvh1o/Ju+rHkkjKekkioHrg4eYNcVry
3iATIJ2ZSdG7I2tMrv+o8Eu7poArUXfJIOL0JRen90VlBEin/petBev2t5n2pkfCRZgN1s0kBFdR
rnyZo87sa+8NiK7IAph+01aHP/upjkjsQ5sOtzdR57AVDm1YhPNNZ6xqrrwwF45/zNKtoNMzTgGP
mwdJsPBapbLI7KYR96eCAsv7wshssTJRVFXsZ+vyYLMZvbPlj+KTFxklQCg7XiswFqcGGq5Fv/oG
u0Rgg86jkrVmbJKZzK8ED90dimFLc8+OHkyUM8q5yX1fgiUkUjw2Olnt0QZq0LXV1QYqScg6jT4l
XozvAQ6tXND/m4axpSypBS9uINkRYap9PcGERb2ifyn35W5gDCypUAU0SUjzUKjb+dZSFMov3934
aCmq8TmwIBRTDLBtjx86vCi4JPQb/4j1V2Z+YzWC9e7aiE0n3ykYsRHiYLNoc1t0BctKVYladmT2
VqsYQb1UWNe5BtrpXtqJWfNcke5/MO4qGRJSEZlyjIaM6A5B0mSboQLJWRWYcSEhw9YUETqx0X3M
E6+FFDF9qaBpZ9ReX5cg+d1Z15YkBw5gB3+fNdfGAs3KmdisjQm18wWZP6dpKEE8FLoA6UC2zybd
sY2I0dr9kMpkT5kQsGWQaJE0ot7Fo6pkoQQDUs+4L1EkGBlTW665wyHVcULJ+QTl6wFA2SBPy8Ee
FD5YmZ+VSZl8i2d9tY3XuZ7mlNDqmBPuwHqT+tD7SDRj79sENBqNmbp4GpjGqbgdbnb2x6ytt2ix
b7SCck+E34IQ/+I5I0voOpGp/H/tb3JS4Byg9TwTmxgdIKePZV0zbYGDIkqoz4veYEJV9Xvj37GH
5GuogRZiHTIqKBaQg2Zs3XKDssz0XspXuofORp3H2PYw5/O+TC394QC2XkjhEy6wnFdXVPPjEOP5
mGtTh3QWBsMzTmWXXG8d7t6bz9RLhFe6+lWSIby7YO2RgmdFf6qi1x8d+biqt3pJvn0aMklN/WHE
XlsIK8gZtiyfVYgm++ZWG/kpXAiI0tQZnjMT2joPqiGz5H/DvwgPGEOo9mnL69HtQZ/xTXJx3yiJ
OnczgaMtZxkNMRz3ZbtTKRgCJ/BOZnxr1MfKMt8crPmizXcVmoYj5KBs0BIgsL7PuFwkQEJPQmrx
eeBADYHwqLhuJGN6TcESxm5YS3fcW4lHyZU3ZuZSqLhKJr9l+4B0B30oWG26tQundfiefZw4HmQW
Y4CYFCvQUX1XV0pfdDK/aY9u5hdekCU/QDECuoXQ6b160KRSoJn6eHWRMDYwJy1gvX+oOT7Czycc
EvZiM+/U1DyryfdGLmS9qVhoCLUbV9qcUYlefj+5I3tcB467HjS5q0wJ5o6YA2N9KklAQ2d24B/B
MVvi3qE2yxkSWIJ5NSrO7P5EQHP/jDz4YJciTa5ZoPdAj9wuY0y5Q4iuFcui4A8Yt1Vw/79BDEo8
yChU3H3us0Rm8/S3XQksyhgNNfUTtyDR9lU2jX4VN/I6sEdlwdNlkVAhwCklBsWDlWKfcxD19UBq
rxo3wZPSRNC2iDbS2iRBX3Pw+55e5SS4AnIMqnnMSggvoOZOycMoYClKyTpxxcDqFZ0TmIhVGz/T
eIolc4ku58bkxA3lnJKN/s+FZfrXNCw6muobTU+nsxcOsTqXYdsVFvoAGOpuCXu3ZE32vbtobLBy
EDrH7WvpurTzI2v7n+4jeA12uUHykWIOZ6o1hLxY3o9j3tPjcDbiKdRJ7m92jOSJONN8s6bXps76
cOQ+OTr+zc+rAKMNdPC3bUYWijxzrgwwd7S9Jp/TZ5fGGhhOdeKwq2Q8iu0KxOX/xQDwpWs3Vi5l
zP5SMaiv9zTzkPASk0+1r1s0bcbYPYgDN+G+ipicsxE5o0PwzS96fVp4Mtun78DO5wTWQQCT5iB5
YcDl4qKiJao3p7mbtWfk0i3zAGyqJz9JdH+VeUTDLv/QVqhks7QcrdJ3KSwsHtXbXkE/FAO7oZHI
tH6ySN5Nn1G9j762ga4wOpZL3npP70fjvf6rOydaMrUrhQAiYwPAUruz5wCBogZiRq7O5cYCsFS9
IwoToelIt7E+6TrOrFfc2RO06cVtrKLcOKgOoMMEsqsZOPDpdk6xqJBsM8BJOokheZ8Axg8c7Ox0
dRkTSZt5Iau9vd2mTFIBuWZbOJefZMDhPxKlAu10CLA/s+px2DYegxRyo4vRnkeDg/24MwrHc++I
PrXTTn2L39lepXKOMi9UvzgM4RKwrdsw7NnyHKD9PR69QLc+IUYD4Po0WPf3S3+hwz5Q4zc8zvgo
/lUbp9M08yTp5duA7pbbNBXQWYgDQxqBasx4VOPSRyn76JfU0nkOuv8CJxp8pnwNoBjBGARy/8La
UNIbZVXvLs6kFxLW4GN+d38GA3S9wGlCNwCZZBBij4gay+0MkRP3qVubrz2Kj3m8bxHJSjT8ELO2
5csPxy4RyGGFExu2osrqL1TsLBQGB/l3313sCBKXnN/3sakOScxZ8UKKAqdAvHnwhLM9RoMkOp5Z
osjChWO1i1STWNaw+1DDVh7/H+Q2CVCuJcaeZo33xBRJVrThdyTUSEXVS5y9HXL86lhNZ5G9MTME
pXtWFye8TM8UdjU+Uq/Edzf8g+5e77eIG2Zt6hzzAFGhllNyZgFALsUT/d5ZIT2ghHtnwOvzWqva
jCFiOnUWhFOzmWrpNSPXDV4Uz+zHhUyVXnb0xRX1R53DKw5HMJfeN0ysHGd12mJeZoRxv9tMcHUn
/NViSXu4Mn7BraYAqrSuU/e/F64iWtqZC6N0XR8XeoD4NB3nRy7LnxxFVXb9wMlOS2QAi+knRSDl
yXxEji6sn0WFIjOP7OGG1prcDUnUI5UW/B9H/TL/1Ikt6ahwIytvKcZ0FEAbHtHCsij5+STOOcY5
+z6ElQIOxWlfHYWED8yhPeZHeAeT3En6TFeRwhmNJvQInhcIhCQVdgnPyp7tkUqEcqQXh9ydbFdM
r4oe9mLyh/qZWOXo1ONBE9jE8TV+u+qipJOdn12eSYIWhDSgtCiMNc09CAHhR8txrTeAGazk3mkK
shsr/Ey4kSdnu0JLp0JIWbO4p/oLA9HP0JJV24Tp6AgDY0CN9/oPmdZ27NF6Gw/IK1GC0jjMIeXy
hE0jy5kXevZKLOf1cGHRoqW50lUrG+CZe1NijhWRc+jE7+bGcATtV5bZNQm5eKYZ6roeChdYL2FA
Gdgge2/6trlWIEVq5zbzyoCN+Nz2VWnS0u8c9xbvovwCfOYYOfH59h3g3kbU+6ufcvh9rDUNokpI
yYRVKeiQL2jNGjvbYbmKB8NcbDOk5rqJ+LTJB6KflkIiyf/I0AK2HdgEaDB/KvWkY6oAEj1uaPlC
KytJTERzRkvz9jYrBxaGT8qi24pqmhdxXa3wMbQakDmmzRwH1BhbO1C31olUC+4yqJfIhBJaFa9D
hmPXaXh4HKH+CEfvBjYPsclX+/rZjdOsVNEs3KT3SrMRqczSgys2W1ls6QsnyjqUCNae98Mquaeo
DoQVqp56x70Dr376pwm4/0OgMIQhcIqc3GiUFsvJTzw/Z5Lb7TB1x96MXWV9bdvWSMOe3EIpl56b
nvgXcOCYDemjnZE1ukOPQ0+f6rkQAemK+GVG4SNlI1/SW5fSCKxXtzcGLxP59tXZ/TfM22bIpbj7
aWTLC0P7Nr7HAPifDyb0j2Wywd1VJkkuETjoDLxqB2gcm2Kd+DnK84IjU3CLSUyJXd1R/ZeWNgne
/12JUw48GDfb8ys6XQGFOUcUj85IkVbcXEQzudHdsj/oQgs6w68i71+AIEYNMZzutONCU6M5m6eW
qDIiYHtnXFe5VdR9wZHOAc2CGHOhuBhaspcyJardv9wbKSbBp4mCphYOVYZ23+7jglEAZYnqdsAO
H5aN0tO07gBUjDdSMdYlzT2MbyA03DgKnP8MT8DBowzEqorlacJtUbSdczSgXmqC5fNpwht9yiPv
XPbnRXKkIR7fGXWCGffZsakFjQUsrGcrBqRgQXVzcsUZ8Wcb0AfBgfQ1JmiFGaTBRcPUQ361geNJ
Kn20+WhvQIqLpx+AiYW+yI1I3Jt6YbiiDtQYS2d7nFdQOJFx0oL4tvmo6HcmqQyYrpg9rmLSJg/0
ErgiHS1txmcLjVphQSu3psc6ROcGfKNJHquebucu8MeeknOPyaVPCqEl5j4aCPAgdJQQjxzdqWGc
zk05qx39wcu/fivv9g7O5k6VuBS8G5FjYWqZPAnNUm1A19WHrp2uCdaZdnM6KCwJVxC+JlaQKfyK
Ad8Xiec7KnLbwDl0SdEaY0O2eXi5fWEmgcoHB8FPDMFLWGhnRwkhdNZEYi58Q8/UDsORP6LdfUh7
AfqFjl8ZrgNQzP7z0vN1WTavGZ4eD5632mh57XuFl0pxE8sk5l7uPWqJPtCeN8YVfkC5bdM/WSSO
LYCoxm6UXJK7l2YYLPeBr3qknTxkU5C5bIqm5xcFxw9rzmZpKvQgE5zcSNyqvO0c6mA9UeWq9280
ZyeQS68CviMdIn5JTP3TpSb5d/Q75/dweg8rEHek52Jzjloec7fAawaRtG+X20KpSO1U4DVAxry8
m1DqmjIVg44B7jn+90JyJeiXh0Yb4oGqDBM+NMrSjLo32C8a4+VMsdVjbICbghZA+k+B6JTJJHsC
zzj2el72/UCAizCtdxEfChU6+pgNZSXWAIfydps3ZW4gvSxrJAXfeMtqX+GMCJodhWXzADpViLLc
gWEb2NyOdYV71SvuZ5akgMfwEA2uMrmhlvLKEb9xSpv7WaxVOwEBGlNXTZhkUZPBQ3Tha25YPfpA
X/l39ccqA6PkHH9O4VyIadshZsQCjfoAD24zoYEacchoX6YpHRkW5foXxguZ52zUEWx9jD4ewysp
V67uXevdyB1pXiYNssYh2cuRY3b2pR/F82QyddsuvQ7U1M8zLc0M5qMRWjbcMkpYHBOEGkyoY1w8
Uo7FTBizM1EaIKjqjXq41VH6bGDfFTQXmeo4uLU7lpW8tn7yU4OBDa73B567Wlqs7evkzaBlj9Ph
MJQQoKQcmPKQYTmPiHF0CzefVyvDmXLB0rQgB+t9oleA0Q6LlRqLk0x6lmRxFa5OkmzdU4Y4c26+
Oo3S52kORkyruw8M8aslHzTUOdSR8QveXMxQKC4ydUi3WuLp7UQbUJTE/GQjkwaH9O26sXOjuKAe
izejBw36cy7ITDmaUqeOMFJ4pRquHdl+vrb81t8X6Ij/aYB91bPaWQ1JXxC71GxwIZ3iDOexAt8B
npAWbN+3bFW3Zd2hiShD3SzHJfnjBmERUi+6V9pPKWscwRsFbO3snMXh3sG+VW2/TK0xdGpKddZQ
JPPzvUuLguA9NmbVsTJlxy/99Qqpe9uoKii2XgQqKkoiuyNXZRmoQ2ePIURsPJQqtKkjnF/KwStn
8NqO6yMGsBWNoJyNOwgaHgQDHoyLV+RvFaYaBw1vRR9N6AP3sclgulPtmFyVlrUuyha/Tq3RxRVE
AoPUpkN9fmykzxlu2l2wjVZv2mqV4jVhKzgmR5YUU5OIvnFU9GONunf36uREZV+ziKwVX2dAJcak
6cSazWKh+65gY00e6m9toLfbUDVXfWKmaMS4hzmVEWovGFGgPYuVBezbO/DHaJcqJPSzC70kLqRw
otEvu3i4vEa3Jg+hIHW6ZeHBdR1uieWrwlXFV8OuA8v/BDCyZP5hhiRD+/sg5LDGbwGPyfbEbqAb
H/5roKOzu5L8UZUi4kwc/xjk3zM31/mSA9d1e/kICR4tzSnRyhNYEC7vNPKR9LTqDjstevbsfwzR
XH8DCP73yOOYFgPRrsiU6+okFWCySK6SWMP1iQ/WEhgUhfx7LfiM8lCpJCE2zTf8GtDos4VhDEye
z36VQDN5jZ548NSqXXS8C+5tAx56H8Gh/pYlGuoQwlxV5tFN3VRK61nxevNxLXvvBxSs3xJL64FL
5xmTtDYPxrhgMIRuIdc51i927s3sJ+buuir0z9KlSI/wrqPXEiTgI4m9gVBBkRI6Jbhw2aS96fcg
ete7lcBB48gypb5BJW3hOpNIdqugCtjy3KHBQR/RXFyxb2N3rFxM57aIZdOLDuzWVSbAK6jq9bm2
4ROBybq70jS7GRW7NHAimvbjOY/Q1ub4h3Agc0k7smngrctpiCpSg1zZTTMx2QetOuuvuRo6PGRD
xz0bdRrdhGWksb+IzdNbLO7oILQ+izl/UdPlhduj8YkcP8b5N3hrws+u6Ket+wjye4qGQfNWNAvW
dfLiwQZmRJD2tExNb5/TsirzBqSxXL77wwCkgl7hM53hCx0/CwrrF2nLE5cuhxzlXSNDh6iwVMcf
9G2MK9aapwpBCphm/hDgHdb8M5tuQxnibShCQ5Cr2sJtetT7w13CEtb5lXeuvxinbeDVhiWywq37
3EhenWzLDf8fSMx7l/Bn5J3aYEoX/o3bUpcnmdAR3QuytGXUxL31yfpL/zBX2lfrLReTa5tRjnIS
V9NuIBXXjThdpGl9eTWEd1fNvUKRzBhn2kdDsV+st7XAbNilZPApLYeFH2xPw6r3+sb+mIrR2Jzu
LJInGr2q4WFMfFbZsTLqXhjZeuT1sK4nCylpCsLN+oDyc23va61+zGLVPEyJN3yBEb87EpHG124B
YqOiOqEYt8doCIxA+ioezTMeX9GOG69zBEYHm7eZvtaL1YqKVxFL8XfWx62sCB4uI8/HYi2awcK5
CuU7f4OmsOOLCA70788ANKHpt36xxgQSBUz4lkVpAfSIZaeE3lGk7W/ZN7INKNG9OAbTjIqfEKEf
X+N/XENtzfSGPxmmiQfJEukjcTUcewgQ4+CrXZFvriJHZwkTsqHgs/DxFz1+pOmuj2DYYEcLu/iI
pZB7bgNMc+z3YGDgZN50WKRBMQzGOXoAK+Gw3OLA3aidlqJkdOGtMKKHWmtI1IXxO8G5I+kuWoNR
4C9wzI3qABcZN2DAhWN/wjN4hqRYUc5SG5g/tm1g1E4BKIzoHLF/N3DlqHTAassNuCsUTU91CjOP
zGTbO18gtmFQPHTi4EBJg+oU2p5hw17GmS338Lk7soqip1uCoRLtgk39phLwKlUYcXZUXaavmxy0
+bFb9PKEIByULFxanjvd1ZgP0xuCMXGnuP6/sxJOlUD/j1vzaLgw/6BeYvCljF0dypbcGrWNji+h
YQDXBZ3SWbVIvZQ5zkkgrhBstFer7OGYbP5djd6VBQFFBMxHkooC1n85Wn4KdSuKg27RfREafViz
/68FNyEyxq3ejTzoUpHkEsJgegoDmnSi9x2u4BWQ27NkEsAXphsA+yWESkl8G/5kO91WgIAxS6PQ
fLOyCCnGP5LsT9HAEhW95NllCRRWmrGFfAu8F+gQJm+ZJ9znQILoHfvY9wG0dG+oavLxCSB9TOAD
+SoGDPluFb+rnxi/Ub5CKUvGCj5MCZgW7CTo5ADLOXfCWfY7j9N5p6TGTTYiYNwAVxKMrZKWsE8i
0qRkqi7WyKmy/GQxu9Q1V9lejHz1PoKHkrTWxBtY/e3Nz+DSSdLA2C5Gqsyx9Wy/zqrVyrnQ7DgM
6uF7PCjh97rpzLlOG60D+OHhKxuaJ2T8RZ97lCF1dAPQstnKMIbXCiX8WEVasF5nMYsTq8WrJ5ff
DsertV7mdRyudh4IF/Yj7VYDXDBSwvCgY1C8pGtalchaL8JzF+T54kq869rMDqezJNlOAqVlP7jd
v63450QSHTDqy3osn203FRb7/x1w1YzbzgVj/5dKGqTnpuzVrmQe74joAhDHP4voAWqa+GdQJAac
fTXu2zZLao4xlDlbWUBz5X4i+5O9Af41J61H/tH1tL5acDuci8DrHecLEeoy05xNfbRsmbmHFjaP
Y1mjWsw0Sc4sWYBrL8YNYhmGGGZW5DFGUX01/A+YVjh4+XgtDNfbeZqoIwYJ/WAFOUBjFjvMMAUw
j2hklkxuuN2a1qPO/Fpd97M3bkNicB5BXEZlsh0N5SgxZAuAFeVxyfxNQVUbOI+paHhA0pDJzVMJ
gsslBy6eBjXrUw605YUtmi1HSYNn/U+tRFAGvraX16b0Tzdu2Gz+ocv6MFXuTcrVw+iwMe00jL5u
XN2HLi4t9blyMyOabvP/2g8rgtERba4Tn6A6ersPDVFVp8VLVpbWBPXcUj6+2jc+CneguWMZFUoc
hTjJL42WBqYAPfLxPLcF6mBBTsaeCEu35lp9Y92lsrWLelqRhTyNZHqC6zDiCcrhPt6SSalZSLzQ
8ivY8OFUI9DhobnboaEYUV1qjGALZP/0XMpYdqDsa+S5jEy4fJ1nFzN2LdYOv1iNZAHndt87GQoq
2sNJLqcjLdfEo6VDfcSlx7Qarqnd6UQv2imLxjLJgtz5wQE6EBnJ1wSwwgUETj4Kst+cksibL8PJ
8+HK58xwSNiPHPtyoFhLFPkq0wIDfs+xDThj/K7vJpApbFvsLUcgZI9FUIj08pday2lIf3L4GR3C
kdb1OVjRSTeOsiBomMjImKP3d6Z4K9YVmr/K8+eO0xc2zThR4hoJWTDzbKCQ0kN+22eqAtlnYtGK
njb5IjwLSwuKwC4Z4mHlpSUSJ7tGZgm6LDnUcmkj44VvdLX2jrSgPpGbpV2maSPPu/JJuBhFYlat
HhzA7u4lMW6QYw4h/iyZPUGk+oVLFA+t2eURcHB4M44TrLZL2JesjBDcSbjW5aUrwQ4Zu+/zV+aX
fX8C5cXY82QH41Kl5pyrA4TSVfTkxRgyCvIr5ZBHrvbyMZPj+UhUC11pVupZ+voR2JmhwXCvpFW3
a3gpoC4GiVxRnejrY9F8bE0xHF+WAESNxuo2+XH7xGZKU62X2XLK4Lh1w+on1Q290FqTXEA6vGIA
hKkN/ad2/rOZx1Mu10JmUI6JzdiO9tOyL92EWhXOt2Qs34PTHtZNrsoI8V6n1Z4nYBjxGN1JmoZc
HEcwiPPy4i6Ywmccm8Nm2oNKahCjjJlxWAEq8E1DVQw9+E3M123/1vubb48HbAfwZFi0nnARw+n5
8INM5/5oEzPLgjXAQO7wAwvM9YQGTjAiIDGRnWpYzb8QmiKiNf4o3oLwQxGRn2B7ZmqX6+n3nedv
3wnAOBksIkWdunGwyNxYuUMxZljMZw/3zvMehau2VPKLGwS0/WTWzoe1mtCzxKnwxwV3Kg5GcWe6
/qxbbrmeOvhi1Aw3+3uatDhDUogJSXlR13SZKAiVliCmMTyBUDfN1//gfN/2x9zTpUs3+M+uODZQ
atxqUlTtrp/55JhFXUaKTSEjkWf8iBD9BtaTkFA4eovERbgDVRburSIdw3yESGu3b/q/IeiAu7Ef
augOOosWHwxDj9ZAaRzXzR+hEJQj1TCh99eStFYT0so9m86EcHjQhqsXAf5K8Gfdp21joc2a+avS
zof0+HUm8cLlYZYo2mSIR2MrlOTujnNS6GjcUf9VqdwGHQRkUryh4IJ3MVMaB0X22S6diLnfcafY
ZZWiudhQ5bzM8fgCbuxB8laZwYI53dqyj1tHnCF/LylYb236szpMix1C3B2fX0xK/VEagy8DNbB4
GWGB+0xB7w2rk++QspAbQVvCXw52sXe3U17/LL+Hal3VqgA2ICuTd0QMWR0pgVja0JjM2mACGeKN
aZB1T+hcl5MHVSv6gDULMZLWuUXnMjGEOy2aHJnNPFKPoc4w3oQJW2oad12N3sauOj0IYZBxREFQ
/zwv2m3X86zcLueGtpsNCoCsv/wuBM0N9xvzBxaXsMf4Q0t643u30GKhmDIgmaHJAaZqtgqFIe/l
hr0jCwqQMKFHAPr6RBeC3Vgb+2vMLvJpmVIyalDK9EsMsHopKuDRT0qLqmBCc0ytH89eiYOveT6Q
SQN2s8yQCiLflCX5rdspAiUS9Vmt9c3969nvTmO7QZqb4lfLGR0/OZqUCph0uFhCTBulvn162jeh
QOJW54yPJVyVfbuykv95l53a13qLW4XKDvlNBI9zsvVPCrrMAzfabdni0X2od2WfsfvaQkz8CPND
TcNT5LS7yy3W/brGuCyFxL8scN3QNtYLaqcYe9w6LSe+5mABetu/v0Yu2SrGKvtEOGni7FkU9AZp
8jef4IevRJKKzUaO4/FFQC3RwSTK4YWRueHAhFbrnRKM3AZPS0uOmyLx+Y9+B6R5YjMZCIrFlCo4
XWOu5EOKPGlwVK5dVhipeoiqTcEPYf3/WIqENCFpxYpf128WLShRY70yh+wtiEZ5SszahYvqEVfU
+bllNm917C5z10So2FQrlaGCwrlg+1/OEf7WkX5zlaeMl3iZ3AICmDNk+zY4KYoOmrOBKNBC5jea
eZmv3JHk/Dp5sTWGFMaK9NfIre1ni+OgxtVBF9YXEJ/i2XM6C388ALcnpsIigAP03Kxwz3tgA6LK
CMQ7YU/Hg+rKQY3k6OqsjAVXBPAAW/YE5gsZFddrIBTDv8B9VxCnbwlvRkBPC14V0ql/oFzI4Gd3
MOr4XN/Sw4oh/vtMOdSNlTACQeKXYGcaVivIc7zaIcFkjADFSgr6ZJsD3m5Uxfys2LEaj7qriwcQ
sxCA6W+h9GXP/YX+h5taJ4zKn01WoQcpH7gVxw1+VX5XPD01qlq0eIv70RtWmrH5mLToory3l+Es
o1mnORNyerzIFhn9pSxN3q1j+a77uYVQUpR79pt1tgy7c2LhXKZueOv338KkdWq4gYcxHkyCYHuf
f0yqKdpbHg8iUzhspjAlkkala28FYzraGURqrNDzVYXdE0V7nDZ7x9bcEyxeFwwCaxSDE6Gsypmd
HkwyWDRsfgbfpUJxv5oKAsNPOsfUBk42xCn1tmEEktBlFF/CSO0wuxfOc2h0NYO2kgOT0i3Xut0c
M1rz6glYT5EnQYuG7CaTGI3F7SDtoK8YmaIYNRrnws4VgRdBBqJhkZAtz5zExZBSyMOa9yoP3w5I
dtaxqtMCIhk1BsWswyvTOwys8fcH6V+H3C3jZSWWAyQLyeLK7jMTHTekwViS3NxNNmullh2Vta8x
IiOQK0AF6AxXI3BQ4mqVCTt3+WgIHQAXxJjv5+1zEhBKtNcOBJBJEFfgGVygPFlS8a8ggKJ1nAL7
LZoVwP2dPhBImsHe6r58MMvfHYBhqTImzGu5TxH3xx8CEAgA5SSsJV5EjFLzy39AC46vu6Jznswy
2GaYcZvgYQqBi/Dda04NfYFPkDWqkwqBdUZIch8iQjcLslK0tPYbd2EKv8MscL4R6Fm/+WEMDJcg
kVkDSx/1/sM6fTeq+kd/3VxP6N+9oy3vi3I8MthcMi6o38hoT74x4j3MZYmiMHOgKfgtEKPNIkL7
DwSCkFrFkNmCME94C43KnWf578LAdEnV2dOWP3ZKXWQnj6OFPU4fy1kE07DEeVzysJgcKPXLK5H+
mkQbSC1ll8+pn6KCc0G9awR6tH0jROj00pbwtVdl6FRqbsLk/jzxCFhJUbjafqf5QnBlvgcEDJB7
t55VzAkcqIRYsdhEL+SKh7Sv0odSthbT19WU2argB+jYVsHjz+Ycwk2a8ar3fdOiqijEc3R0Xh2N
sEq/3nCW9x0G6/dP3pnfplxCgogH7+Wdgv4C7v+7yrEh8MG8q31RecHyWckN+jc5VT3YAt45Clb/
2b2U6vns9VAqC1UdvJiw2BP7EQtea+MofJAxgxlD2ACKWfl/e5H6aIpZl2W6jgn0NSOU8maQ3Dsb
WFBn4OdYjvDDiCyDO0lVmWVhihg3YndamWi4mvEY9fy8BwSGeu1vr3KNEoxr84m85r/E1xxKdXYN
lFhnI7sN83DWBO9Z55MFtgoVoMgKIrmA5piaZi+WHnrt2KFSfrQbJJxa5AsEbdITh9UY6DVhIZ3g
PSArQpcGQtssZHcgt7UgLNOQVxEmcjUfmKHDOhkb2HNlhMuw/pxGk0lWyRENqe6gqzc6ObEqKggA
U+2RnDuJM85l22G88sRbPI5b1mlDwTP20O7a1f/M510v4WkqQqb98cxduyFX2OUdpFfr5crQBrpC
TxeOXApW6YbGoeejN4d27dLBHg92mPC/oK9IPexRU4FKCDBKkhNjn2YhcCsfavXZ+koAyKWS+tOU
IbIK5djfdYAIrCHNPe0SiiFEFUNhJ7QjktQIPGLtT6pwi65tiobMYoH5d7Jnw004XhicdUd4FGnS
EwhZkzi7GF+47pCLJIFsiz6071gP8h432FwRLmrp4V5oIR3MtJV9Qwo0aLD2qu0KKZ4mkdK+k5KI
j3DTPz5gWFZ/2bWSY6do+JdsP6gp037SHYN5FyxfO+BnrGjYRtlQPBiM8ssvcjDvDXr+XzR6OGjX
puZVaS8RPiBBl2dPfAlXy9JAA/xFtRYRtYjQLn7ybm68gRgSidXacTMW+dHsbYXKYE+hsqaHYQps
JvGEsOKSTS6RZfZbIcAKKeC2oJmZk0fAQ546CpRXYwrN8OgHxvO/gl9NfOGFs5l1B5+OhLuPnlzg
x3aADsY0QI3XeVpX6flNtPFgJ3EmmdWeq2R5XUVBSxKpNtdBPNppY0VHFpjyuVw2wZLB4tyzCSy4
XhV2d4I4cpKtH6OR7dC6h8prxqBulmgEKupiRbHjtc5Ek9uVnbSoawezz3sgLbp8x8NpaTwFwdI0
2vDQQw9quGuE3h0sdaz8U7WKXHGnh3KyUkBDxFsIhGR++/qUoQU8kkVtusBYwsIhivHEASrPT/0/
o03r4KPteDTxdBoCIsn4xadGsxsfDDZaarilw4/4+cqMK7H3StIl2gFZC7+JEYpLxCrRVscS8Si+
b4qdCcPIUQZQqn41uwR2AsIz/ynLaIgrUwam8RIxOuJqdsw0/2aUQdgaKHRs/vz2p/zlvK+zcxMt
5ibVSqW/xBw9FlORgIsImJWXgsrtgowoK0PwZR5CznZ8w5XX4HqlUX2zmqOED64Tlgls7d70IfSM
AQBIYJqZ26T9d4aln8Z2eIRpToRVB1EMOAuuZzEKmsP0bXTDnRu55Gsjvn3SCQmA5ABHyjFOVeGQ
U4Zr9iuqxcrm6evddmjSQBjpGxqBSe4A/Eh1BjSR3Cpp4F1RgVSyBvx0MrFUSTlCkOZ9TF4t9Gbj
rN/J8ThO8X6ssQPMIiFn/twyZ0Q09j0UD1WatbPbOn4GIMByhHlmikNWpmaZ/Rr+7Csa+ehPhQta
w3tSJnxTT+hc8AMETC1BlIn6aO7lkevey5B58hQJ8W/OeCoHEsRsLFyM5EZ5DYVC5KuqEZNCI9Qh
ByEi+Wgow47VPgt+vNxp3edaF2Fzeft85aSNTbyuzmtC8NUXTGt7vqY4D0azIvh3X3WRDmpnD/L8
tfwX90EuVllVaQxQIPwVqwaRVBeAmQgrOWVhBv5AwMFYsXP8fReRaExdjVq4htEU6fpN7Z1dYQBI
/O3Ko5fnJPLX0AHq68fD5kCixu8heS09sTMLeMQvkdXusPafPYUNUQeU1no4xI8a6zLtDrWD+wX/
ULEjL3pBlDWUmr8zJvupQTnvh1LazHytD4KrxPfc1DSQKmGSbTqLnv2j7w9FTsxhArkOaM9hKnYE
8KLxeBp/KJb0Ol2k2KVhXWNh7RBzilqVCKu52kIXNR06Nqf2jptTTMU6AnVnhu38XIfLjVCV2d5T
cO0frktzGh1/t8D0ah3fP0VBU+A7HxHjR1y9b69n9JV6vTFVp2jhhtPdorZV2y4NM8+ZTd7ExTAz
KvaTZCQLMBaEhi7biXLjCxqyhB7/Mq++hECU/QEIT+iiJFOLyfwtw9tJoeFL/zLOkXjyEhZdOdrY
NF4TrCRtPCCZCjOT9uqWTOFL/K4mxG6NFA1f2sJomhmAzlngKj+z/+Z7W4hsY8FPfLkUrVLAsei9
1fEq45plNRKwzCU6yIuGZd1W3JdlgxcSm6425H8LFYGXsqTczXd4Obwa3M2kw7TRkt/QgSBWX8Dm
6ooI7/5OaW1XgXBPVwG6CncqN/KwjysfT3xNx+RtSk49LTtOKb3JroUw/X7nWZMXJzmC1YcCeruu
YcNq5wTWJZT53lOjVAD/8S5kz3NMPkUazVSrey9clQXnj4gWiYKHropnUyuTL2funTx/MxMF+5hg
ZOaeUepoNN1xpSrCaYHow11/e2TuKQu0G/2JLwzwR91LK7Jss2a5zn7QX+AEsIcaP4wefqUjiJq6
tZIAJqfxXX8ziWLn8wsh6T70BcIPijHBtH5R91dpD5cU+MAt5c6ZJ1EYHhoGzskl8NxEUkypuFxb
5oWrp7pZ/NvfUWEpViV6QPF2a+Tn5aWZiFTnCl0GYyve57dQ8nf4F22DMxuygobHMIwiYYqbXxV/
II/Uq0jPCFpvOU7nSDuf2OTs3rsoULaZAnmyYASvOmFyEH27wFA7dK1mGB54SOY7W/gl55eVs2Kj
NhyG/8/MN9le9KjZHxadmnZjYVtB/IVVMLJ4Cfk6uf3+v/im/huQdoIzqAm/2ja8QBxuiJcwsIxT
kCwziCaT/kxPP6NkW89xmE7OzYA70mM3+CsY49zRB4U5nRu0TDykBo/vxkVe9tJAO5cIS8Yf5nB3
eQrvfKA0dSzH+1ArNZpjeWk3mNDLHRVNPcnJbIy9FSLhVoyA4YIHy0LqyJq0WKjPRGQ1mASEDOiI
whfdjIHlPLJfdWFTKo9PhjDQr+mpZiHUZH1C3niNgBcxhYOcxkeYL6tnwEHv7eQLXmK/vwJRZOJy
rIpsuDVSpihX8YxpZRG/f5LfY/j88sJpv6EOEjBwNJRKEwqIIyEkFFurvIU8vsdnmaavOgrhiFyP
FwvFPPAJiGvSxg5s4loBxo7jrfkD/v3o0wufv+mqXn/wSpJA9iWTDXKd79LmZj/IsAuI31wIWGpy
B7BDNn7/DwC6sIEo/1fpoBqkL1O22UVzonhg9+VjERw4O581GRlAeeAEfgvmOUW6igrRN/kFb7V2
eUR1DVIxb+syqzOoWCBph14CmePP/hTP/eCYA1U7B7WYKEf22/ydAbMhOGjEYSDDDyMuZiZtjf1C
vBZfjHzRSBKgrhcpkeBe+nxJUKRfErGi8oc06vjo2eS7fc1rzF2+GzqHEASms+7QjnuCa63/jGNn
htN28ruIJjBqMnVcljkHLf7EI0L+W+leWWe6xK+PFgJcvlm+M30bETsnoR9W41kPL0t+cbiJWiKR
m62fixe5ck96lcBMiEBAxtzdqNKSbPjHOOxYyb1szmjaz0HDs5jKlEnH2ajPd1wOzqz2eKNE+w/T
mxVXtw4/I32lRQ8uKUHcV3wL6t3Z0vAh/fnNN13WJQB24rGjhTi97Vw8ON2TSC7/4PIhsD057FVZ
trlEsqbwt74SKSFPun75V8wmZlC7IvQGSViDrfFkenO4vbx9KTa2i+Op/KNeZ5SejqHmNRYlRCdC
DlF4AG9ycDldY86AsgRAVRlrT7bKrYgI1k0TkUTwSInIlG1fJkJbybNdIXKUhQHThkamVRbna8tL
jEbwbgSpuk2oxgr2K3enWVFq5PNe6nIrgUtRmZ2mVQByzjTmTyVjCatSD5l6gsS3oIbialL3smFm
lX2yHMzv1sGuCfjwKCuhVHrcxYsdbkcxfW5GsvnL+ZjgzzTvByrUcqtZ83zZm8KMxhI4iAONVeh7
OAZYNBPhK5PksNT9ebHdWKO35eKbp5WVYwVYIP5UGGXLUFrpJj08ed+oRRdRDfDjKlxc36ETQTvG
4hoEf7iV4b59aifiK0lPTF0CsLmzao+b0i5IwuljnxEgyqwXWWcayzNf/m41qRpY185FWZ76hKfL
UKBjpxYsha7I68gmDQREoPvzf8s9kA8T6UzhbsPsj+wGnDo+bHlCwoKUiDXE8q6+Z3W2m+eqVBbS
+AnxX9MOtDBPRhc+IyDqLN5SZIKzULDQQgbhEsAvX9XVf4EZ4Wxsr6BSCWBGdpj7Pl63H7IwroGE
xvqQ2PGIjN56DnRTHXqxkgWLc42WcpQpekY90lK/b6NzuZs8mjUGZnd83sRQe/734HH7PKEOxoca
Q/D4XPEXggMVlnIy3AmXBjv3PFv9r3pp7233lP1iNWtwuAU8L/3HXjufRDg+GpSe7NGPfStz5/aV
uTlOg19PZp49sZF9uB9wl0mDHJdDgXXVHE1mnHgZWGxap1R1i2eCz1uou6cfXOJ8MIYVb15T4udA
auyu2JVCkb10DiBKH3UqWRLpfK4CS29c6I5mVYpV7Skw4NrKEVEcKyEAB8PKWp+ImQyum4pFN6wz
4gfc1jZSjMf+lQQ2b9CJhtk45F9cf94c/f2py3Blhzz5naXYZ5bbj5wZS0ltBRZ0sE9OQ5ZnBtrZ
ypfqoV1E7ahabJ8/eYbuRsmoDhHJxq7You63yu7NKgUAMF4vaADcGh9lWqJANJgAJ1naT5Pn8V8V
jBpGnSxSDYIaT0aUv6m0gP33lmdCWKnqUmKfLd6ot2ClnPNne9OjT6ZLbsGOGbAJg2hekzDg4mLJ
XCvZNnTDZ42aiH0qG8XVGIk+qtv7wopeszJiacHKGQUhuqO3HvReNsd/I5/HL5HjT3S5w8vwGM6M
RfBXtM3IKqOpjH4DS/qooW065/zzAb/8krwMTY5RYkMLbWZD6CRDtUkvRNWrwBLAtJkEb6vwHfs2
5pNlD1ooRmG4EFv/fPvl8QWxXwHHR50WtVrdDXQQsMR4FbY2Axu+ImdzwRtCNtM9liO53dI972B9
bj+JHSz0Q/1lt4Nrk+HRtsi4PkzqqgHXjqXLe7rXeL/5BfhGSxZxMPFU7jxbulsXvco6we/5Pqqb
rInDoLHMOV8U1LN/U0T6dblOdz3yKDjGdevlStcZQe3XKL9EpG+LjlZgUEOUwLZhTxrmbVBdgR75
aCmKR98LRm0NHIkPe0Iw1u4NJixAYQ8qcy/Q9Pog+aJddr1tfkCg3y3EdNSVyslVmk6FD2jMJXFM
AAhTQc8jmHLg9+he671Jh1gWdgZ5Lpagbf6bTvOUsAvUnLcGr/L7viiKUdCXZ9Z8sNPJxd9kyPfE
/auOyZePVn3XHtRmUM/IIOBNzKX7z8vVwRxzX6OAyXHMkn7LDSd5xQ/voykQxN6koUVWdAuDCl7A
wpdvy5g/Ksoxa3bMjt+Nn3gJAIlPLn+Ntv+Qxz4r5hgE4/tdD4OPyS7S4HKXX3UmEP6prIuGdjng
tci27AFpuzI+ziMpzD/zlfJnbcXqZcW0qCLg8ngwwixe0fljqGk7DrDi0BEXALkvT0TQLJNb+P5f
nkbhEevH13v7A7qhNaVH9dIeSNAsiPTG0zEd9UI7XK1UOSYBuOJfFH9MY5oQxox2z4ViWnO3Agxd
kE6RFnsmtuOEx7C2QUSJ6MxDMBFp3NH3ZFsPJpr87vIMqWkImVvx4q+yUcl07kUT/2ZRqNDkJxDk
XqM347X/jBhIdlttPXdEMsV2tqf9sp3N6o4khTvTjHYttheoDQhliSYezluO3H3PgluFYGDWCuIx
9RElgaI9Bu6+4BOK0lbfCMuzonlpfoia+278utSjWM1QqG8crbdR1GTktfccDEGEeWG/lg+B7Crt
7el5LL3JJkvry//AiH+N1ceWNzQbwFy/XvO3CyvmygMNEhxdQkfg8lBfQtpd0ZCZSHx6FD5gjy8j
U18qSi7aBtVig48I//mgA2BbqcD6NLq06PKcaQEqm+Zau/6cqy8AobWRgD9Ix+pEDSztkST6qXdI
34YoX0FI/3PnWgIOS9C9EgeXqHbvLLEQcih5QxtOw+XOAIM0W+7z8G235eRau/PyIkyAR8G28WsO
wilZPqwuSojzPlEmXEVpalY00t3ydBgI8Zaxoc0NF6TA4EUOHtfjvUAKhpWyr58cpWJzEIGnFt95
lt5sABaCZ0TskD/ccS8nB6OJklyKBWbKnWiuAN6E4E1Kzbjq0+r5OG/8X8431rWofAqgkpxJ4Cqn
WFQUrOSl98DCwkKmYIVeFRu5kQNXBnQIheeIlm+9OgBhvnA5PD/4913fsxegWuvRC715tU+C85/E
vSY7waT6DEyd4esc5ESvOt1oUPnkbexFa5qOkJxjWS/kAJwcBqdiuBFGd+QT7lSbt5f7CemTEvWY
d4tGnhECLt0TG8IUZwPzm36XuIIwy/NlCb0JuH8zNCtl3fg=
`pragma protect end_protected
